`timescale 10ns / 1ns

//purely combinational array of multiplexers
module interconnect #(parameter WIDTH =4) (
input wire [31:0] control_signal,                 // 2-bit control signal to select Weight/Input stationary as well as Uni/Multicast modes
input wire [ WIDTH-1:0] stationary_signal_1,     // 81 Weight/Input stationary signal that will be broadcasted to all PE's
input wire [ WIDTH-1:0] stationary_signal_2,
input wire [ WIDTH-1:0] stationary_signal_3,
input wire [ WIDTH-1:0] stationary_signal_4,
input wire [ WIDTH-1:0] stationary_signal_5,
input wire [ WIDTH-1:0] stationary_signal_6,
input wire [ WIDTH-1:0] stationary_signal_7,
input wire [ WIDTH-1:0] stationary_signal_8,
input wire [ WIDTH-1:0] stationary_signal_9,
input wire [ WIDTH-1:0] stationary_signal_10,
input wire [ WIDTH-1:0] stationary_signal_11,
input wire [ WIDTH-1:0] stationary_signal_12,
input wire [ WIDTH-1:0] stationary_signal_13,
input wire [ WIDTH-1:0] stationary_signal_14,
input wire [ WIDTH-1:0] stationary_signal_15,
input wire [ WIDTH-1:0] stationary_signal_16,
input wire [ WIDTH-1:0] stationary_signal_17,
input wire [ WIDTH-1:0] stationary_signal_18,
input wire [ WIDTH-1:0] stationary_signal_19,
input wire [ WIDTH-1:0] stationary_signal_20,
input wire [ WIDTH-1:0] stationary_signal_21,
input wire [ WIDTH-1:0] stationary_signal_22,
input wire [ WIDTH-1:0] stationary_signal_23,
input wire [ WIDTH-1:0] stationary_signal_24,
input wire [ WIDTH-1:0] stationary_signal_25,
input wire [ WIDTH-1:0] stationary_signal_26,
input wire [ WIDTH-1:0] stationary_signal_27,
input wire [ WIDTH-1:0] stationary_signal_28,
input wire [ WIDTH-1:0] stationary_signal_29,
input wire [ WIDTH-1:0] stationary_signal_30,
input wire [ WIDTH-1:0] stationary_signal_31,
input wire [ WIDTH-1:0] stationary_signal_32,
input wire [ WIDTH-1:0] stationary_signal_33,
input wire [ WIDTH-1:0] stationary_signal_34,
input wire [ WIDTH-1:0] stationary_signal_35,
input wire [ WIDTH-1:0] stationary_signal_36,
input wire [ WIDTH-1:0] stationary_signal_37,
input wire [ WIDTH-1:0] stationary_signal_38,
input wire [ WIDTH-1:0] stationary_signal_39,
input wire [ WIDTH-1:0] stationary_signal_40,
input wire [ WIDTH-1:0] stationary_signal_41,
input wire [ WIDTH-1:0] stationary_signal_42,
input wire [ WIDTH-1:0] stationary_signal_43,
input wire [ WIDTH-1:0] stationary_signal_44,
input wire [ WIDTH-1:0] stationary_signal_45,
input wire [ WIDTH-1:0] stationary_signal_46,
input wire [ WIDTH-1:0] stationary_signal_47,
input wire [ WIDTH-1:0] stationary_signal_48,
input wire [ WIDTH-1:0] stationary_signal_49,
input wire [ WIDTH-1:0] stationary_signal_50,
input wire [ WIDTH-1:0] stationary_signal_51,
input wire [ WIDTH-1:0] stationary_signal_52,
input wire [ WIDTH-1:0] stationary_signal_53,
input wire [ WIDTH-1:0] stationary_signal_54,
input wire [ WIDTH-1:0] stationary_signal_55,
input wire [ WIDTH-1:0] stationary_signal_56,
input wire [ WIDTH-1:0] stationary_signal_57,
input wire [ WIDTH-1:0] stationary_signal_58,
input wire [ WIDTH-1:0] stationary_signal_59,
input wire [ WIDTH-1:0] stationary_signal_60,
input wire [ WIDTH-1:0] stationary_signal_61,
input wire [ WIDTH-1:0] stationary_signal_62,
input wire [ WIDTH-1:0] stationary_signal_63,
input wire [ WIDTH-1:0] stationary_signal_64,
input wire [ WIDTH-1:0] stationary_signal_65,          
input wire [ WIDTH-1:0] stationary_signal_66,
input wire [ WIDTH-1:0] stationary_signal_67,
input wire [ WIDTH-1:0] stationary_signal_68,
input wire [ WIDTH-1:0] stationary_signal_69,
input wire [ WIDTH-1:0] stationary_signal_70,
input wire [ WIDTH-1:0] stationary_signal_71,
input wire [ WIDTH-1:0] stationary_signal_72,
input wire [ WIDTH-1:0] stationary_signal_73,
input wire [ WIDTH-1:0] stationary_signal_74,
input wire [ WIDTH-1:0] stationary_signal_75,
input wire [ WIDTH-1:0] stationary_signal_76,
input wire [ WIDTH-1:0] stationary_signal_77,
input wire [ WIDTH-1:0] stationary_signal_78,
input wire [ WIDTH-1:0] stationary_signal_79,
input wire [ WIDTH-1:0] stationary_signal_80,
input wire [ WIDTH-1:0] stationary_signal_81,
input wire [ WIDTH-1:0] sw_input_1,              // 81 Weight/Input  signals that will be uni/multicasted to all PE's
input wire [ WIDTH-1:0] sw_input_2,
input wire [ WIDTH-1:0] sw_input_3,
input wire [ WIDTH-1:0] sw_input_4,
input wire [ WIDTH-1:0] sw_input_5,
input wire [ WIDTH-1:0] sw_input_6,
input wire [ WIDTH-1:0] sw_input_7,
input wire [ WIDTH-1:0] sw_input_8,
input wire [ WIDTH-1:0] sw_input_9,
input wire [ WIDTH-1:0] sw_input_10,
input wire [ WIDTH-1:0] sw_input_11,
input wire [ WIDTH-1:0] sw_input_12,
input wire [ WIDTH-1:0] sw_input_13,
input wire [ WIDTH-1:0] sw_input_14,
input wire [ WIDTH-1:0] sw_input_15,
input wire [ WIDTH-1:0] sw_input_16,
input wire [ WIDTH-1:0] sw_input_17,
input wire [ WIDTH-1:0] sw_input_18,
input wire [ WIDTH-1:0] sw_input_19,
input wire [ WIDTH-1:0] sw_input_20,
input wire [ WIDTH-1:0] sw_input_21,
input wire [ WIDTH-1:0] sw_input_22,
input wire [ WIDTH-1:0] sw_input_23,
input wire [ WIDTH-1:0] sw_input_24,
input wire [ WIDTH-1:0] sw_input_25,
input wire [ WIDTH-1:0] sw_input_26,
input wire [ WIDTH-1:0] sw_input_27,
input wire [ WIDTH-1:0] sw_input_28,
input wire [ WIDTH-1:0] sw_input_29,
input wire [ WIDTH-1:0] sw_input_30,
input wire [ WIDTH-1:0] sw_input_31,
input wire [ WIDTH-1:0] sw_input_32,
input wire [ WIDTH-1:0] sw_input_33,
input wire [ WIDTH-1:0] sw_input_34,
input wire [ WIDTH-1:0] sw_input_35,
input wire [ WIDTH-1:0] sw_input_36,
input wire [ WIDTH-1:0] sw_input_37,
input wire [ WIDTH-1:0] sw_input_38,
input wire [ WIDTH-1:0] sw_input_39,
input wire [ WIDTH-1:0] sw_input_40,
input wire [ WIDTH-1:0] sw_input_41,
input wire [ WIDTH-1:0] sw_input_42,
input wire [ WIDTH-1:0] sw_input_43,
input wire [ WIDTH-1:0] sw_input_44,
input wire [ WIDTH-1:0] sw_input_45,
input wire [ WIDTH-1:0] sw_input_46,
input wire [ WIDTH-1:0] sw_input_47,
input wire [ WIDTH-1:0] sw_input_48,
input wire [ WIDTH-1:0] sw_input_49,
input wire [ WIDTH-1:0] sw_input_50,
input wire [ WIDTH-1:0] sw_input_51,
input wire [ WIDTH-1:0] sw_input_52,
input wire [ WIDTH-1:0] sw_input_53,
input wire [ WIDTH-1:0] sw_input_54,
input wire [ WIDTH-1:0] sw_input_55,
input wire [ WIDTH-1:0] sw_input_56,
input wire [ WIDTH-1:0] sw_input_57,
input wire [ WIDTH-1:0] sw_input_58,
input wire [ WIDTH-1:0] sw_input_59,
input wire [ WIDTH-1:0] sw_input_60,
input wire [ WIDTH-1:0] sw_input_61,
input wire [ WIDTH-1:0] sw_input_62,
input wire [ WIDTH-1:0] sw_input_63,
input wire [ WIDTH-1:0] sw_input_64,
input wire [ WIDTH-1:0] sw_input_65,          
input wire [ WIDTH-1:0] sw_input_66,
input wire [ WIDTH-1:0] sw_input_67,
input wire [ WIDTH-1:0] sw_input_68,
input wire [ WIDTH-1:0] sw_input_69,
input wire [ WIDTH-1:0] sw_input_70,
input wire [ WIDTH-1:0] sw_input_71,
input wire [ WIDTH-1:0] sw_input_72,
input wire [ WIDTH-1:0] sw_input_73,
input wire [ WIDTH-1:0] sw_input_74,
input wire [ WIDTH-1:0] sw_input_75,
input wire [ WIDTH-1:0] sw_input_76,
input wire [ WIDTH-1:0] sw_input_77,
input wire [ WIDTH-1:0] sw_input_78,
input wire [ WIDTH-1:0] sw_input_79,
input wire [ WIDTH-1:0] sw_input_80,
input wire [ WIDTH-1:0] sw_input_81,
input wire [6:0] index_1,                 //   81 index signals to select target MAC Unit
input wire [6:0] index_2,
input wire [6:0] index_3,
input wire [6:0] index_4,
input wire [6:0] index_5,
input wire [6:0] index_6,
input wire [6:0] index_7,
input wire [6:0] index_8,
input wire [6:0] index_9,
input wire [6:0] index_10,
input wire [6:0] index_11,
input wire [6:0] index_12,
input wire [6:0] index_13,
input wire [6:0] index_14,
input wire [6:0] index_15,
input wire [6:0] index_16,
input wire [6:0] index_17,
input wire [6:0] index_18,
input wire [6:0] index_19,
input wire [6:0] index_20,
input wire [6:0] index_21,
input wire [6:0] index_22,
input wire [6:0] index_23,
input wire [6:0] index_24,
input wire [6:0] index_25,
input wire [6:0] index_26,
input wire [6:0] index_27,
input wire [6:0] index_28,
input wire [6:0] index_29,
input wire [6:0] index_30,
input wire [6:0] index_31,
input wire [6:0] index_32,
input wire [6:0] index_33,
input wire [6:0] index_34,
input wire [6:0] index_35,
input wire [6:0] index_36,
input wire [6:0] index_37,
input wire [6:0] index_38,
input wire [6:0] index_39,
input wire [6:0] index_40,
input wire [6:0] index_41,
input wire [6:0] index_42,
input wire [6:0] index_43,
input wire [6:0] index_44,
input wire [6:0] index_45,
input wire [6:0] index_46,
input wire [6:0] index_47,
input wire [6:0] index_48,
input wire [6:0] index_49,
input wire [6:0] index_50,
input wire [6:0] index_51,
input wire [6:0] index_52,
input wire [6:0] index_53,
input wire [6:0] index_54,
input wire [6:0] index_55,
input wire [6:0] index_56,
input wire [6:0] index_57,
input wire [6:0] index_58,
input wire [6:0] index_59,
input wire [6:0] index_60,
input wire [6:0] index_61,
input wire [6:0] index_62,
input wire [6:0] index_63,
input wire [6:0] index_64,
input wire [6:0] index_65,
input wire [6:0] index_66,
input wire [6:0] index_67,
input wire [6:0] index_68,
input wire [6:0] index_69,
input wire [6:0] index_70,
input wire [6:0] index_71,
input wire [6:0] index_72,
input wire [6:0] index_73,
input wire [6:0] index_74,
input wire [6:0] index_75,
input wire [6:0] index_76,
input wire [6:0] index_77,
input wire [6:0] index_78,
input wire [6:0] index_79,
input wire [6:0] index_80,
input wire [6:0] index_81,  
output wire [ WIDTH-1:0] sw_output_1,           //   162 output signals from interconnect that goes to the pe_array
output wire [ WIDTH-1:0] sw_output_2,
output wire [ WIDTH-1:0] sw_output_3,
output wire [ WIDTH-1:0] sw_output_4,
output wire [ WIDTH-1:0] sw_output_5,
output wire [ WIDTH-1:0] sw_output_6,
output wire [ WIDTH-1:0] sw_output_7,
output wire [ WIDTH-1:0] sw_output_8,
output wire [ WIDTH-1:0] sw_output_9,
output wire [ WIDTH-1:0] sw_output_10,
output wire [ WIDTH-1:0] sw_output_11,
output wire [ WIDTH-1:0] sw_output_12,
output wire [ WIDTH-1:0] sw_output_13,
output wire [ WIDTH-1:0] sw_output_14,
output wire [ WIDTH-1:0] sw_output_15,
output wire [ WIDTH-1:0] sw_output_16,
output wire [ WIDTH-1:0] sw_output_17,
output wire [ WIDTH-1:0] sw_output_18,
output wire [ WIDTH-1:0] sw_output_19,
output wire [ WIDTH-1:0] sw_output_20,
output wire [ WIDTH-1:0] sw_output_21,
output wire [ WIDTH-1:0] sw_output_22,
output wire [ WIDTH-1:0] sw_output_23,
output wire [ WIDTH-1:0] sw_output_24,
output wire [ WIDTH-1:0] sw_output_25,
output wire [ WIDTH-1:0] sw_output_26,
output wire [ WIDTH-1:0] sw_output_27,
output wire [ WIDTH-1:0] sw_output_28,
output wire [ WIDTH-1:0] sw_output_29,
output wire [ WIDTH-1:0] sw_output_30,
output wire [ WIDTH-1:0] sw_output_31,
output wire [ WIDTH-1:0] sw_output_32,
output wire [ WIDTH-1:0] sw_output_33,
output wire [ WIDTH-1:0] sw_output_34,
output wire [ WIDTH-1:0] sw_output_35,
output wire [ WIDTH-1:0] sw_output_36,
output wire [ WIDTH-1:0] sw_output_37,
output wire [ WIDTH-1:0] sw_output_38,
output wire [ WIDTH-1:0] sw_output_39,
output wire [ WIDTH-1:0] sw_output_40,
output wire [ WIDTH-1:0] sw_output_41,
output wire [ WIDTH-1:0] sw_output_42,
output wire [ WIDTH-1:0] sw_output_43,
output wire [ WIDTH-1:0] sw_output_44,
output wire [ WIDTH-1:0] sw_output_45,
output wire [ WIDTH-1:0] sw_output_46,
output wire [ WIDTH-1:0] sw_output_47,
output wire [ WIDTH-1:0] sw_output_48,
output wire [ WIDTH-1:0] sw_output_49,
output wire [ WIDTH-1:0] sw_output_50,
output wire [ WIDTH-1:0] sw_output_51,
output wire [ WIDTH-1:0] sw_output_52,
output wire [ WIDTH-1:0] sw_output_53,
output wire [ WIDTH-1:0] sw_output_54,
output wire [ WIDTH-1:0] sw_output_55,
output wire [ WIDTH-1:0] sw_output_56,
output wire [ WIDTH-1:0] sw_output_57,
output wire [ WIDTH-1:0] sw_output_58,
output wire [ WIDTH-1:0] sw_output_59,
output wire [ WIDTH-1:0] sw_output_60,
output wire [ WIDTH-1:0] sw_output_61,
output wire [ WIDTH-1:0] sw_output_62,
output wire [ WIDTH-1:0] sw_output_63,
output wire [ WIDTH-1:0] sw_output_64,
output wire [ WIDTH-1:0] sw_output_65,          
output wire [ WIDTH-1:0] sw_output_66,
output wire [ WIDTH-1:0] sw_output_67,
output wire [ WIDTH-1:0] sw_output_68,
output wire [ WIDTH-1:0] sw_output_69,
output wire [ WIDTH-1:0] sw_output_70,
output wire [ WIDTH-1:0] sw_output_71,
output wire [ WIDTH-1:0] sw_output_72,
output wire [ WIDTH-1:0] sw_output_73,
output wire [ WIDTH-1:0] sw_output_74,
output wire [ WIDTH-1:0] sw_output_75,
output wire [ WIDTH-1:0] sw_output_76,
output wire [ WIDTH-1:0] sw_output_77,
output wire [ WIDTH-1:0] sw_output_78,
output wire [ WIDTH-1:0] sw_output_79,
output wire [ WIDTH-1:0] sw_output_80,
output wire [ WIDTH-1:0] sw_output_81,
output wire [ WIDTH-1:0] sw_output_82,
output wire [ WIDTH-1:0] sw_output_83,
output wire [ WIDTH-1:0] sw_output_84,
output wire [ WIDTH-1:0] sw_output_85,
output wire [ WIDTH-1:0] sw_output_86,
output wire [ WIDTH-1:0] sw_output_87,
output wire [ WIDTH-1:0] sw_output_88,
output wire [ WIDTH-1:0] sw_output_89,
output wire [ WIDTH-1:0] sw_output_90,
output wire [ WIDTH-1:0] sw_output_91,
output wire [ WIDTH-1:0] sw_output_92,
output wire [ WIDTH-1:0] sw_output_93,
output wire [ WIDTH-1:0] sw_output_94,
output wire [ WIDTH-1:0] sw_output_95,
output wire [ WIDTH-1:0] sw_output_96,
output wire [ WIDTH-1:0] sw_output_97,
output wire [ WIDTH-1:0] sw_output_98,
output wire [ WIDTH-1:0] sw_output_99,
output wire [ WIDTH-1:0] sw_output_100,
output wire [ WIDTH-1:0] sw_output_101,
output wire [ WIDTH-1:0] sw_output_102,
output wire [ WIDTH-1:0] sw_output_103,
output wire [ WIDTH-1:0] sw_output_104,
output wire [ WIDTH-1:0] sw_output_105,
output wire [ WIDTH-1:0] sw_output_106,
output wire [ WIDTH-1:0] sw_output_107,
output wire [ WIDTH-1:0] sw_output_108,
output wire [ WIDTH-1:0] sw_output_109,
output wire [ WIDTH-1:0] sw_output_110,
output wire [ WIDTH-1:0] sw_output_111,
output wire [ WIDTH-1:0] sw_output_112,
output wire [ WIDTH-1:0] sw_output_113,
output wire [ WIDTH-1:0] sw_output_114,
output wire [ WIDTH-1:0] sw_output_115,
output wire [ WIDTH-1:0] sw_output_116,
output wire [ WIDTH-1:0] sw_output_117,
output wire [ WIDTH-1:0] sw_output_118,
output wire [ WIDTH-1:0] sw_output_119,
output wire [ WIDTH-1:0] sw_output_120,
output wire [ WIDTH-1:0] sw_output_121,
output wire [ WIDTH-1:0] sw_output_122,
output wire [ WIDTH-1:0] sw_output_123,
output wire [ WIDTH-1:0] sw_output_124,
output wire [ WIDTH-1:0] sw_output_125,
output wire [ WIDTH-1:0] sw_output_126,
output wire [ WIDTH-1:0] sw_output_127,
output wire [ WIDTH-1:0] sw_output_128,
output wire [WIDTH-1:0] sw_output_129,
output wire [WIDTH-1:0] sw_output_130,
output wire [WIDTH-1:0] sw_output_131,
output wire [WIDTH-1:0] sw_output_132,
output wire [WIDTH-1:0] sw_output_133,
output wire [WIDTH-1:0] sw_output_134,
output wire [WIDTH-1:0] sw_output_135,
output wire [WIDTH-1:0] sw_output_136,
output wire [WIDTH-1:0] sw_output_137,
output wire [WIDTH-1:0] sw_output_138,
output wire [WIDTH-1:0] sw_output_139,
output wire [WIDTH-1:0] sw_output_140,
output wire [WIDTH-1:0] sw_output_141,
output wire [WIDTH-1:0] sw_output_142,
output wire [WIDTH-1:0] sw_output_143,
output wire [WIDTH-1:0] sw_output_144,
output wire [WIDTH-1:0] sw_output_145,
output wire [WIDTH-1:0] sw_output_146,
output wire [WIDTH-1:0] sw_output_147,
output wire [WIDTH-1:0] sw_output_148,
output wire [WIDTH-1:0] sw_output_149,
output wire [WIDTH-1:0] sw_output_150,
output wire [WIDTH-1:0] sw_output_151,
output wire [WIDTH-1:0] sw_output_152,
output wire [WIDTH-1:0] sw_output_153,
output wire [WIDTH-1:0] sw_output_154,
output wire [WIDTH-1:0] sw_output_155,
output wire [WIDTH-1:0] sw_output_156,
output wire [WIDTH-1:0] sw_output_157,
output wire [WIDTH-1:0] sw_output_158,
output wire [WIDTH-1:0] sw_output_159,
output wire [WIDTH-1:0] sw_output_160,
output wire [WIDTH-1:0] sw_output_161,
output wire [WIDTH-1:0] sw_output_162                   
);
//for the first 81 outputs weights are either broadcasted/unicasted or multicasted 
 assign sw_output_1 =   (control_signal[1] == 0) ? stationary_signal_1:                                     // for weight matrix broadcasting in weight stationary mode
                        (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :                     // for input multi/uni cast in input stationary mode
                        (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                        (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                        (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                        (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                        (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                        (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 : 
                        (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :
                        (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 :
                        
                        (control_signal[0] ==0&& index_1 == 7'b0000001) ? sw_input_1 : 
                        (control_signal[0] ==0&& index_2 == 7'b0000001) ? sw_input_2 : 
                        (control_signal[0] ==0&& index_3 == 7'b0000001) ? sw_input_3 : 
                        (control_signal[0] ==0&& index_4 == 7'b0000001) ? sw_input_4 : 
                        (control_signal[0] ==0&& index_5 == 7'b0000001) ? sw_input_5 : 
                        (control_signal[0] ==0&& index_6 == 7'b0000001) ? sw_input_6 : 
                        (control_signal[0] ==0&& index_7 == 7'b0000001) ? sw_input_7 : 
                        (control_signal[0] ==0&& index_8 == 7'b0000001) ? sw_input_8 :              
                        (control_signal[0] ==0&& index_9 == 7'b0000001) ? sw_input_9 : 
                        (control_signal[0] ==0&& index_10 == 7'b0000001) ? sw_input_10 : 
                        (control_signal[0] ==0&& index_11 == 7'b0000001) ? sw_input_11 : 
                        (control_signal[0] ==0&& index_12 == 7'b0000001) ? sw_input_12 : 
                        (control_signal[0] ==0&& index_13 == 7'b0000001) ? sw_input_13 : 
                        (control_signal[0] ==0&& index_14 == 7'b0000001) ? sw_input_14 : 
                        (control_signal[0] ==0&& index_15 == 7'b0000001) ? sw_input_15 : 
                        (control_signal[0] ==0&& index_16 == 7'b0000001) ? sw_input_16 : 
                        (control_signal[0] ==0&& index_17 == 7'b0000001) ? sw_input_17: 
                        (control_signal[0] ==0&& index_18 == 7'b0000001) ? sw_input_18 : 
                        (control_signal[0] ==0&& index_19 == 7'b0000001) ? sw_input_19 : 
                        (control_signal[0] ==0&& index_20 == 7'b0000001) ? sw_input_20 : 
                        (control_signal[0] ==0&& index_21 == 7'b0000001) ? sw_input_21 : 
                        (control_signal[0] ==0&& index_22 == 7'b0000001) ? sw_input_22 : 
                        (control_signal[0] ==0&& index_23 == 7'b0000001) ? sw_input_23 : 
                        (control_signal[0] ==0&& index_24 == 7'b0000001) ? sw_input_24 : 
                        (control_signal[0] ==0&& index_25 == 7'b0000001) ? sw_input_25 : 
                        (control_signal[0] ==0&& index_26 == 7'b0000001) ? sw_input_26 : 
                        (control_signal[0] ==0&& index_27 == 7'b0000001) ? sw_input_27 : 
                        (control_signal[0] ==0&& index_28 == 7'b0000001) ? sw_input_28 : 
                        (control_signal[0] ==0&& index_29 == 7'b0000001) ? sw_input_29 : 
                        (control_signal[0] ==0&& index_30 == 7'b0000001) ? sw_input_30 : 
                        (control_signal[0] ==0&& index_31 == 7'b0000001) ? sw_input_31 : 
                        (control_signal[0] ==0&& index_32 == 7'b0000001) ? sw_input_32 : 
                        (control_signal[0] ==0&& index_33 == 7'b0000001) ? sw_input_33 : 
                        (control_signal[0] ==0&& index_34 == 7'b0000001) ? sw_input_34 : 
                        (control_signal[0] ==0&& index_35 == 7'b0000001) ? sw_input_35 : 
                        (control_signal[0] ==0&& index_36 == 7'b0000001) ? sw_input_36 : 
                        (control_signal[0] ==0&& index_37 == 7'b0000001) ? sw_input_37 : 
                        (control_signal[0] ==0&& index_38 == 7'b0000001) ? sw_input_38 : 
                        (control_signal[0] ==0&& index_39 == 7'b0000001) ? sw_input_39 : 
                        (control_signal[0] ==0&& index_40 == 7'b0000001) ? sw_input_40 : 
                        (control_signal[0] ==0&& index_41 == 7'b0000001) ? sw_input_41 : 
                        (control_signal[0] ==0&& index_42 == 7'b0000001) ? sw_input_42 : 
                        (control_signal[0] ==0&& index_43 == 7'b0000001) ? sw_input_43 : 
                        (control_signal[0] ==0&& index_44 == 7'b0000001) ? sw_input_44 : 
                        (control_signal[0] ==0&& index_45 == 7'b0000001) ? sw_input_45 : 
                        (control_signal[0] ==0&& index_46 == 7'b0000001) ? sw_input_46 : 
                        (control_signal[0] ==0&& index_47 == 7'b0000001) ? sw_input_47 : 
                        (control_signal[0] ==0&& index_48 == 7'b0000001) ? sw_input_48 : 
                        (control_signal[0] ==0&& index_49 == 7'b0000001) ? sw_input_49 : 
                        (control_signal[0] ==0&& index_50 == 7'b0000001) ? sw_input_50 : 
                        (control_signal[0] ==0&& index_51 == 7'b0000001) ? sw_input_51 : 
                        (control_signal[0] ==0&& index_52 == 7'b0000001) ? sw_input_52 : 
                        (control_signal[0] ==0&& index_53 == 7'b0000001) ? sw_input_53 : 
                        (control_signal[0] ==0&& index_54 == 7'b0000001) ? sw_input_54 : 
                        (control_signal[0] ==0&& index_55 == 7'b0000001) ? sw_input_55 : 
                        (control_signal[0] ==0&& index_56 == 7'b0000001) ? sw_input_56 : 
                        (control_signal[0] ==0&& index_57 == 7'b0000001) ? sw_input_57 : 
                        (control_signal[0] ==0&& index_58 == 7'b0000001) ? sw_input_58 : 
                        (control_signal[0] ==0&& index_59 == 7'b0000001) ? sw_input_59 : 
                        (control_signal[0] ==0&& index_60 == 7'b0000001) ? sw_input_60 : 
                        (control_signal[0] ==0&& index_61 == 7'b0000001) ? sw_input_61 : 
                        (control_signal[0] ==0&& index_62 == 7'b0000001) ? sw_input_62 : 
                        (control_signal[0] ==0&& index_63 == 7'b0000001) ? sw_input_63 : 
                        (control_signal[0] ==0&& index_64 == 7'b0000001) ? sw_input_64 :   
                        (control_signal[0] ==0&& index_65 == 7'b0000001) ? sw_input_65 : 
                        (control_signal[0] ==0&& index_66 == 7'b0000001) ? sw_input_66 : 
                        (control_signal[0] ==0&& index_67 == 7'b0000001) ? sw_input_67 : 
                        (control_signal[0] ==0&& index_68 == 7'b0000001) ? sw_input_68 : 
                        (control_signal[0] ==0&& index_69 == 7'b0000001) ? sw_input_69 : 
                        (control_signal[0] ==0&& index_70 == 7'b0000001) ? sw_input_70 : 
                        (control_signal[0] ==0&& index_71 == 7'b0000001) ? sw_input_71 : 
                        (control_signal[0] ==0&& index_72 == 7'b0000001) ? sw_input_72 : 
                        (control_signal[0] ==0&& index_73 == 7'b0000001) ? sw_input_73 : 
                        (control_signal[0] ==0&& index_74 == 7'b0000001) ? sw_input_74 : 
                        (control_signal[0] ==0&& index_75 == 7'b0000001) ? sw_input_75 : 
                        (control_signal[0] ==0&& index_76 == 7'b0000001) ? sw_input_76 : 
                        (control_signal[0] ==0&& index_77 == 7'b0000001) ? sw_input_77 : 
                        (control_signal[0] ==0&& index_78 == 7'b0000001) ? sw_input_78 :  
                        (control_signal[0] ==0&& index_79 == 7'b0000001) ? sw_input_79 : 
                        (control_signal[0] ==0&& index_80 == 7'b0000001) ? sw_input_80 : 
                        (control_signal[0] ==0&& index_81 == 7'b0000001) ? sw_input_81 :            
                        7'bzzzzzzz; 
assign sw_output_2 =    (control_signal[1] == 0) ? stationary_signal_2:               
                        (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                        (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                        (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                        (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                        (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                        (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                        (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 : 
                        (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :
                        (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 :
                        
                        (control_signal[0] ==0&& index_1 == 7'b0000010) ? sw_input_1 : 
                        (control_signal[0] ==0&& index_2 == 7'b0000010) ? sw_input_2 : 
                        (control_signal[0] ==0&& index_3 == 7'b0000010) ? sw_input_3 : 
                        (control_signal[0] ==0&& index_4 == 7'b0000010) ? sw_input_4 : 
                        (control_signal[0] ==0&& index_5 == 7'b0000010) ? sw_input_5 : 
                        (control_signal[0] ==0&& index_6 == 7'b0000010) ? sw_input_6 : 
                        (control_signal[0] ==0&& index_7 == 7'b0000010) ? sw_input_7 : 
                        (control_signal[0] ==0&& index_8 == 7'b0000010) ? sw_input_8 :              
                        (control_signal[0] ==0&& index_9 == 7'b0000010) ? sw_input_9 : 
                        (control_signal[0] ==0&& index_10 == 7'b0000010) ? sw_input_10 : 
                        (control_signal[0] ==0&& index_11 == 7'b0000010) ? sw_input_11 : 
                        (control_signal[0] ==0&& index_12 == 7'b0000010) ? sw_input_12 : 
                        (control_signal[0] ==0&& index_13 == 7'b0000010) ? sw_input_13 : 
                        (control_signal[0] ==0&& index_14 == 7'b0000010) ? sw_input_14 : 
                        (control_signal[0] ==0&& index_15 == 7'b0000010) ? sw_input_15 : 
                        (control_signal[0] ==0&& index_16 == 7'b0000010) ? sw_input_16 : 
                        (control_signal[0] ==0&& index_17 == 7'b0000010) ? sw_input_17: 
                        (control_signal[0] ==0&& index_18 == 7'b0000010) ? sw_input_18 : 
                        (control_signal[0] ==0&& index_19 == 7'b0000010) ? sw_input_19 : 
                        (control_signal[0] ==0&& index_20 == 7'b0000010) ? sw_input_20 : 
                        (control_signal[0] ==0&& index_21 == 7'b0000010) ? sw_input_21 : 
                        (control_signal[0] ==0&& index_22 == 7'b0000010) ? sw_input_22 : 
                        (control_signal[0] ==0&& index_23 == 7'b0000010) ? sw_input_23 : 
                        (control_signal[0] ==0&& index_24 == 7'b0000010) ? sw_input_24 : 
                        (control_signal[0] ==0&& index_25 == 7'b0000010) ? sw_input_25 : 
                        (control_signal[0] ==0&& index_26 == 7'b0000010) ? sw_input_26 : 
                        (control_signal[0] ==0&& index_27 == 7'b0000010) ? sw_input_27 : 
                        (control_signal[0] ==0&& index_28 == 7'b0000010) ? sw_input_28 : 
                        (control_signal[0] ==0&& index_29 == 7'b0000010) ? sw_input_29 : 
                        (control_signal[0] ==0&& index_30 == 7'b0000010) ? sw_input_30 : 
                        (control_signal[0] ==0&& index_31 == 7'b0000010) ? sw_input_31 : 
                        (control_signal[0] ==0&& index_32 == 7'b0000010) ? sw_input_32 : 
                        (control_signal[0] ==0&& index_33 == 7'b0000010) ? sw_input_33 : 
                        (control_signal[0] ==0&& index_34 == 7'b0000010) ? sw_input_34 : 
                        (control_signal[0] ==0&& index_35 == 7'b0000010) ? sw_input_35 : 
                        (control_signal[0] ==0&& index_36 == 7'b0000010) ? sw_input_36 : 
                        (control_signal[0] ==0&& index_37 == 7'b0000010) ? sw_input_37 : 
                        (control_signal[0] ==0&& index_38 == 7'b0000010) ? sw_input_38 : 
                        (control_signal[0] ==0&& index_39 == 7'b0000010) ? sw_input_39 : 
                        (control_signal[0] ==0&& index_40 == 7'b0000010) ? sw_input_40 : 
                        (control_signal[0] ==0&& index_41 == 7'b0000010) ? sw_input_41 : 
                        (control_signal[0] ==0&& index_42 == 7'b0000010) ? sw_input_42 : 
                        (control_signal[0] ==0&& index_43 == 7'b0000010) ? sw_input_43 : 
                        (control_signal[0] ==0&& index_44 == 7'b0000010) ? sw_input_44 : 
                        (control_signal[0] ==0&& index_45 == 7'b0000010) ? sw_input_45 : 
                        (control_signal[0] ==0&& index_46 == 7'b0000010) ? sw_input_46 : 
                        (control_signal[0] ==0&& index_47 == 7'b0000010) ? sw_input_47 : 
                        (control_signal[0] ==0&& index_48 == 7'b0000010) ? sw_input_48 : 
                        (control_signal[0] ==0&& index_49 == 7'b0000010) ? sw_input_49 : 
                        (control_signal[0] ==0&& index_50 == 7'b0000010) ? sw_input_50 : 
                        (control_signal[0] ==0&& index_51 == 7'b0000010) ? sw_input_51 : 
                        (control_signal[0] ==0&& index_52 == 7'b0000010) ? sw_input_52 : 
                        (control_signal[0] ==0&& index_53 == 7'b0000010) ? sw_input_53 : 
                        (control_signal[0] ==0&& index_54 == 7'b0000010) ? sw_input_54 : 
                        (control_signal[0] ==0&& index_55 == 7'b0000010) ? sw_input_55 : 
                        (control_signal[0] ==0&& index_56 == 7'b0000010) ? sw_input_56 : 
                        (control_signal[0] ==0&& index_57 == 7'b0000010) ? sw_input_57 : 
                        (control_signal[0] ==0&& index_58 == 7'b0000010) ? sw_input_58 : 
                        (control_signal[0] ==0&& index_59 == 7'b0000010) ? sw_input_59 : 
                        (control_signal[0] ==0&& index_60 == 7'b0000010) ? sw_input_60 : 
                        (control_signal[0] ==0&& index_61 == 7'b0000010) ? sw_input_61 : 
                        (control_signal[0] ==0&& index_62 == 7'b0000010) ? sw_input_62 : 
                        (control_signal[0] ==0&& index_63 == 7'b0000010) ? sw_input_63 : 
                        (control_signal[0] ==0&& index_64 == 7'b0000010) ? sw_input_64 : 
                        (control_signal[0] ==0&& index_65 == 7'b0000010) ? sw_input_65 : 
                        (control_signal[0] ==0&& index_66 == 7'b0000010) ? sw_input_66 : 
                        (control_signal[0] ==0&& index_67 == 7'b0000010) ? sw_input_67 : 
                        (control_signal[0] ==0&& index_68 == 7'b0000010) ? sw_input_68 : 
                        (control_signal[0] ==0&& index_69 == 7'b0000010) ? sw_input_69 : 
                        (control_signal[0] ==0&& index_70 == 7'b0000010) ? sw_input_70 : 
                        (control_signal[0] ==0&& index_71 == 7'b0000010) ? sw_input_71 : 
                        (control_signal[0] ==0&& index_72 == 7'b0000010) ? sw_input_72 : 
                        (control_signal[0] ==0&& index_73 == 7'b0000010) ? sw_input_73 : 
                        (control_signal[0] ==0&& index_74 == 7'b0000010) ? sw_input_74 : 
                        (control_signal[0] ==0&& index_75 == 7'b0000010) ? sw_input_75 : 
                        (control_signal[0] ==0&& index_76 == 7'b0000010) ? sw_input_76 : 
                        (control_signal[0] ==0&& index_77 == 7'b0000010) ? sw_input_77 : 
                        (control_signal[0] ==0&& index_78 == 7'b0000010) ? sw_input_78 :  
                        (control_signal[0] ==0&& index_79 == 7'b0000010) ? sw_input_79 : 
                        (control_signal[0] ==0&& index_80 == 7'b0000010) ? sw_input_80 : 
                        (control_signal[0] ==0&& index_81 == 7'b0000010) ? sw_input_81 :                                                 
                         7'bzzzzzzz; 
assign sw_output_3 =  (control_signal[1] == 0) ? stationary_signal_3:              
                      (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0000011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0000011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0000011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0000011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0000011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0000011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0000011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0000011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0000011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0000011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0000011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0000011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0000011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0000011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0000011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0000011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0000011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0000011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0000011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0000011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0000011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0000011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0000011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0000011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0000011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0000011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0000011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0000011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0000011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0000011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0000011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0000011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0000011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0000011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0000011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0000011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0000011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0000011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0000011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0000011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0000011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0000011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0000011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0000011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0000011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0000011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0000011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0000011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0000011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0000011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0000011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0000011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0000011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0000011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0000011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0000011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0000011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0000011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0000011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0000011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0000011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0000011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0000011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0000011) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0000011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0000011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0000011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0000011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0000011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0000011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0000011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0000011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0000011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0000011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0000011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0000011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0000011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0000011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0000011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0000011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0000011) ? sw_input_81 :                                  
                      7'bzzzzzzz; 
assign sw_output_4 =(control_signal[1] == 0) ? stationary_signal_4:                   
                    (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                    (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                    (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                    (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                    (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                    (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                    (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 : 
                    (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :
                    (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0000100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0000100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0000100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0000100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0000100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0000100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0000100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0000100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0000100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0000100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0000100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0000100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0000100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0000100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0000100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0000100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0000100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0000100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0000100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0000100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0000100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0000100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0000100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0000100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0000100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0000100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0000100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0000100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0000100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0000100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0000100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0000100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0000100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0000100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0000100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0000100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0000100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0000100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0000100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0000100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0000100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0000100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0000100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0000100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0000100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0000100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0000100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0000100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0000100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0000100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0000100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0000100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0000100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0000100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0000100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0000100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0000100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0000100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0000100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0000100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0000100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0000100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0000100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0000100) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0000100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0000100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0000100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0000100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0000100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0000100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0000100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0000100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0000100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0000100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0000100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0000100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0000100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0000100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0000100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0000100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0000100) ? sw_input_81 :                     
                      7'bzzzzzzz;  
assign sw_output_5 =(control_signal[1] == 0) ? stationary_signal_5:
                    (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                    (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                    (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                    (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                    (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                    (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                    (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 : 
                    (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :
                    (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0000101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0000101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0000101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0000101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0000101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0000101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0000101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0000101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0000101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0000101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0000101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0000101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0000101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0000101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0000101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0000101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0000101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0000101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0000101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0000101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0000101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0000101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0000101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0000101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0000101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0000101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0000101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0000101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0000101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0000101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0000101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0000101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0000101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0000101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0000101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0000101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0000101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0000101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0000101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0000101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0000101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0000101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0000101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0000101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0000101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0000101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0000101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0000101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0000101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0000101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0000101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0000101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0000101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0000101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0000101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0000101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0000101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0000101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0000101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0000101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0000101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0000101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0000101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0000101) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0000101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0000101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0000101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0000101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0000101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0000101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0000101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0000101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0000101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0000101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0000101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0000101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0000101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0000101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0000101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0000101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0000101) ? sw_input_81 :                        
                    7'bzzzzzzz; 
assign sw_output_6 =(control_signal[1] == 0) ? stationary_signal_6:                
                    (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                    (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                    (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                    (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                    (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                    (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                    (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 : 
                    (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :
                    (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0000110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0000110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0000110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0000110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0000110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0000110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0000110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0000110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0000110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0000110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0000110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0000110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0000110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0000110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0000110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0000110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0000110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0000110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0000110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0000110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0000110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0000110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0000110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0000110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0000110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0000110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0000110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0000110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0000110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0000110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0000110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0000110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0000110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0000110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0000110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0000110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0000110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0000110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0000110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0000110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0000110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0000110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0000110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0000110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0000110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0000110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0000110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0000110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0000110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0000110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0000110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0000110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0000110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0000110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0000110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0000110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0000110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0000110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0000110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0000110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0000110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0000110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0000110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0000110) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0000110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0000110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0000110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0000110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0000110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0000110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0000110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0000110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0000110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0000110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0000110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0000110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0000110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0000110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0000110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0000110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0000110) ? sw_input_81 :                                                  
                      7'bzzzzzzz;   
assign sw_output_7 =(control_signal[1] == 0) ? stationary_signal_7:                 
                    (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1:
                    (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                    (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                    (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                    (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                    (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                    (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 : 
                    (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :
                    (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0000111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0000111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0000111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0000111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0000111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0000111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0000111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0000111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0000111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0000111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0000111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0000111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0000111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0000111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0000111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0000111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0000111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0000111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0000111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0000111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0000111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0000111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0000111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0000111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0000111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0000111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0000111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0000111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0000111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0000111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0000111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0000111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0000111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0000111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0000111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0000111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0000111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0000111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0000111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0000111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0000111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0000111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0000111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0000111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0000111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0000111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0000111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0000111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0000111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0000111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0000111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0000111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0000111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0000111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0000111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0000111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0000111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0000111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0000111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0000111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0000111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0000111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0000111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0000111) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0000111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0000111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0000111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0000111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0000111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0000111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0000111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0000111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0000111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0000111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0000111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0000111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0000111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0000111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0000111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0000111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0000111) ? sw_input_81 :                           
                     7'bzzzzzzz; 
assign sw_output_8 =  (control_signal[1] == 0) ? stationary_signal_8:                   
                      (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 :
                       
                    (control_signal[0] ==0&& index_1 == 7'b0001000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001000) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0001000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001000) ? sw_input_81 :                              
                      7'bzzzzzzz; 
assign sw_output_9 =  (control_signal[1] == 0) ? stationary_signal_9:                  
                      (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001001) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0001001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001001) ? sw_input_81 :   
                      7'bzzzzzzz; 
assign sw_output_10 = (control_signal[1] == 0) ? stationary_signal_1:                     
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001010) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0001010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001010) ? sw_input_81 :
                      7'bzzzzzzz;   
assign sw_output_11 = (control_signal[1] == 0) ? stationary_signal_2:                  
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001011) ? sw_input_64 : 
                     (control_signal[0] ==0&& index_65 == 7'b0001011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001011) ? sw_input_81 :                                           
                      7'bzzzzzzz; 
assign sw_output_12 = (control_signal[1] == 0) ? stationary_signal_3:                 
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001100) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0001100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001100) ? sw_input_81 : 
                    7'bzzzzzzz;                         
assign sw_output_13 = (control_signal[1] == 0) ? stationary_signal_4:                      
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001101) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0001101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001101) ? sw_input_81 :                      
                    7'bzzzzzzz; 
assign sw_output_14 = (control_signal[1] == 0) ? stationary_signal_5:                       
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001110) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0001110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001110) ? sw_input_81 :                       
                    7'bzzzzzzz; 
assign sw_output_15 = (control_signal[1] == 0) ? stationary_signal_6:                 
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001111) ? sw_input_64 :
                      (control_signal[0] ==0&& index_65 == 7'b0001111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001111) ? sw_input_81 : 
                    7'bzzzzzzz; 
assign sw_output_16 = (control_signal[1] == 0) ? stationary_signal_7:                    
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0010000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010000) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0010000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010000) ? sw_input_81 :                     
                    7'bzzzzzzz;   
assign sw_output_17 = (control_signal[1] == 0) ? stationary_signal_8:
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0010001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010001) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0010001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010001) ? sw_input_81 :                                             
                    7'bzzzzzzz; 
assign sw_output_18 = (control_signal[1] == 0) ? stationary_signal_9: 
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 :   
                      
                    (control_signal[0] ==0&& index_1 == 7'b0010010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010010) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0010010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010010) ? sw_input_81 : 
                    7'bzzzzzzz;                       
assign sw_output_19 = (control_signal[1] == 0) ? stationary_signal_1:
                      (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0010011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010011) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0010011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010011) ? sw_input_81 :                     
                     7'bzzzzzzz; 
assign sw_output_20 = (control_signal[1] == 0) ? stationary_signal_2:
                      (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0010100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010100) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0010100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010100) ? sw_input_81 :               
                    7'bzzzzzzz; 
assign sw_output_21 = (control_signal[1] == 0) ? stationary_signal_3:
                      (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0010101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010101) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0010101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010101) ? sw_input_81 : 
                    7'bzzzzzzz; 
assign sw_output_22 = (control_signal[1] == 0) ? stationary_signal_4:
                      (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0010110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010110) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0010110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010110) ? sw_input_81 :                                           
                    7'bzzzzzzz;   
assign sw_output_23 = (control_signal[1] == 0) ? stationary_signal_5:
                      (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0010111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010111) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0010111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010111) ? sw_input_81 :                       
                    7'bzzzzzzz; 
assign sw_output_24 = (control_signal[1] == 0) ? stationary_signal_6:
                      (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0011000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011000) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0011000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011000) ? sw_input_81 :                     
                    7'bzzzzzzz;                         
assign sw_output_25 = (control_signal[1] == 0) ? stationary_signal_7:
                      (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0011001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011001) ? sw_input_64 : 
                     (control_signal[0] ==0&& index_65 == 7'b0011001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011001) ? sw_input_81 :                                              
                    7'bzzzzzzz; 
assign sw_output_26 = (control_signal[1] == 0) ? stationary_signal_8:
                      (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0011010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011010) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0011010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011010) ? sw_input_81 :              
                    7'bzzzzzzz; 
assign sw_output_27 = (control_signal[1] == 0) ? stationary_signal_9:
                      (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0011011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011011) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0011011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011011) ? sw_input_81 :
                    7'bzzzzzzz; 
assign sw_output_28 = (control_signal[1] == 0) ? stationary_signal_1:
                      (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0011100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011100) ? sw_input_64 :
                     (control_signal[0] ==0&& index_65 == 7'b0011100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011100) ? sw_input_81 :                 
                    7'bzzzzzzz;   
assign sw_output_29 = (control_signal[1] == 0) ? stationary_signal_2:
                      (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0011101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011101) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0011101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011101) ? sw_input_81 :                   
                    7'bzzzzzzz; 
assign sw_output_30 = (control_signal[1] == 0) ? stationary_signal_3:
                      (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0011110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011110) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0011110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011110) ? sw_input_81 :                                            
                     7'bzzzzzzz;                         
assign sw_output_31 = (control_signal[1] == 0) ? stationary_signal_4:
                      (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0011111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011111) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0011111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011111) ? sw_input_81 :                    
                     7'bzzzzzzz; 
assign sw_output_32 = (control_signal[1] == 0) ? stationary_signal_5:
                      (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0100000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100000) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0100000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100000) ? sw_input_81 :          
                    7'bzzzzzzz; 
assign sw_output_33 = (control_signal[1] == 0) ? stationary_signal_6:
                      (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0100001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100001) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100001) ? sw_input_81 :                   
                    7'bzzzzzzz; 
assign sw_output_34 = (control_signal[1] == 0) ? stationary_signal_7:
                      (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0100010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100010) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100010) ? sw_input_81 :             
                     7'bzzzzzzz;   
assign sw_output_35 = (control_signal[1] == 0) ? stationary_signal_8:
                      (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0100011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100011) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100011) ? sw_input_81 :               
                    7'bzzzzzzz; 
assign sw_output_36 = (control_signal[1] == 0) ? stationary_signal_9:
                      (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0100100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100100) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100100) ? sw_input_81 :                 
                    7'bzzzzzzz;                         
assign sw_output_37 = (control_signal[1] == 0) ? stationary_signal_1:
                      (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0100101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100101) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100101) ? sw_input_81 :                      
                     7'bzzzzzzz; 
assign sw_output_38 = (control_signal[1] == 0) ? stationary_signal_2:
                      (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0100110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100110) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100110) ? sw_input_81 :                    
                      7'bzzzzzzz; 
assign sw_output_39 = (control_signal[1] == 0) ? stationary_signal_3:
                      (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0100111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100111) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100111) ? sw_input_81 :
                    7'bzzzzzzz; 
assign sw_output_40 = (control_signal[1] == 0) ? stationary_signal_4:
                      (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0101000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101000) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101000) ? sw_input_81 :               
                    7'bzzzzzzz;   
assign sw_output_41 = (control_signal[1] == 0) ? stationary_signal_5:
                      (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0101001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101001) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101001) ? sw_input_81 :                  
                    7'bzzzzzzz; 
assign sw_output_42 = (control_signal[1] == 0) ? stationary_signal_6:
                      (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0101010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101010) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101010) ? sw_input_81 :               
                    7'bzzzzzzz;                         
assign sw_output_43 = (control_signal[1] == 0) ? stationary_signal_7:
                      (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0101011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101011) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101011) ? sw_input_81 :                 
                    7'bzzzzzzz; 
assign sw_output_44 = (control_signal[1] == 0) ? stationary_signal_8:
                      (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0101100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101100) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101100) ? sw_input_81 :                                           
                    7'bzzzzzzz; 
assign sw_output_45 = (control_signal[1] == 0) ? stationary_signal_9:
                      (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0101101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101101) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101101) ? sw_input_81 : 
                    7'bzzzzzzz; 
assign sw_output_46 = (control_signal[1] == 0) ? stationary_signal_1:
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0101110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101110) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101110) ? sw_input_81 :             
                    7'bzzzzzzz;   
assign sw_output_47 = (control_signal[1] == 0) ? stationary_signal_2:
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0101111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101111) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101111) ? sw_input_81 :             
                    7'bzzzzzzz; 
assign sw_output_48 = (control_signal[1] == 0) ? stationary_signal_3:
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0110000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110000) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110000) ? sw_input_81 :                     
                    7'bzzzzzzz;                         
assign sw_output_49 = (control_signal[1] == 0) ? stationary_signal_4:
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0110001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110001) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110001) ? sw_input_81 :                    
                    7'bzzzzzzz; 
assign sw_output_50 = (control_signal[1] == 0) ? stationary_signal_5:
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0110010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110010) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110010) ? sw_input_81 :                   
                    7'bzzzzzzz; 
assign sw_output_51 = (control_signal[1] == 0) ? stationary_signal_6:
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0110011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110011) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110001) ? sw_input_81 :
                    7'bzzzzzzz; 
assign sw_output_52 = (control_signal[1] == 0) ? stationary_signal_7:
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0110100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110100) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110100) ? sw_input_81 :                
                    7'bzzzzzzz;   
assign sw_output_53 = (control_signal[1] == 0) ? stationary_signal_8:                   
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                      
                      
                    (control_signal[0] ==0&& index_1 == 7'b0110101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110101) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110101) ? sw_input_81 :                  
                    7'bzzzzzzz; 
assign sw_output_54 = (control_signal[1] == 0) ? stationary_signal_9:
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0110110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110110) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110110) ? sw_input_81 :             
                    7'bzzzzzzz;                         
assign sw_output_55 = (control_signal[1] == 0) ? stationary_signal_1:
                      (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0110111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110111) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110111) ? sw_input_81 :                 
                    7'bzzzzzzz; 
assign sw_output_56 = (control_signal[1] == 0) ? stationary_signal_2:                   
                      (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0111000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111000) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0111000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111000) ? sw_input_81 :                      
                    7'bzzzzzzz; 
assign sw_output_57 = (control_signal[1] == 0) ? stationary_signal_3:                  
                      (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                     
                    (control_signal[0] ==0&& index_1 == 7'b0111001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111001) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0111001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111001) ? sw_input_81 :  
                    7'bzzzzzzz; 
assign sw_output_58 = (control_signal[1] == 0) ? stationary_signal_4:                  
                      (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                     
                    (control_signal[0] ==0&& index_1 == 7'b0111010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111010) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0111010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111010) ? sw_input_81 :                     
                    7'bzzzzzzz;   
assign sw_output_59 = (control_signal[1] == 0) ? stationary_signal_5:                  
                      (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0111011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111011) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0111011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111011) ? sw_input_81 :                         
                    7'bzzzzzzz; 
assign sw_output_60 = (control_signal[1] == 0) ? stationary_signal_6:                   
                      (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0111100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111100) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0111100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111100) ? sw_input_81 :                         
                    7'bzzzzzzz;                         
assign sw_output_61 = (control_signal[1] == 0) ? stationary_signal_7:                   
                      (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0111101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111101) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0111101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111101) ? sw_input_81 :                        
                    7'bzzzzzzz; 
assign sw_output_62 = (control_signal[1] == 0) ? stationary_signal_8:              
                      (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0111110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111110) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0111110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111110) ? sw_input_81 :                       
                    7'bzzzzzzz; 
assign sw_output_63 = (control_signal[1] == 0) ? stationary_signal_9:                   
                      (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0111111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111111) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0111111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111111) ? sw_input_81 : 
                     7'bzzzzzzz; 
assign sw_output_64 = (control_signal[1] == 0) ? stationary_signal_1:    
                      (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :  
                      
                    (control_signal[0] ==0&& index_1 == 7'b1000000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1000000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1000000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1000000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1000000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1000000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1000000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1000000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1000000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1000000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1000000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1000000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1000000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1000000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1000000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1000000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1000000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1000000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1000000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1000000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1000000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1000000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1000000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1000000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1000000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1000000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1000000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1000000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1000000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1000000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1000000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1000000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1000000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1000000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1000000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1000000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1000000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1000000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1000000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1000000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1000000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1000000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1000000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1000000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1000000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1000000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1000000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1000000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1000000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1000000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1000000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1000000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1000000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1000000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1000000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1000000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1000000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1000000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1000000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1000000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1000000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1000000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1000000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1000000) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b1000000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1000000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1000000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1000000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1000000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1000000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1000000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1000000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1000000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1000000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1000000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1000000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1000000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1000000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1000000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1000000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000000) ? sw_input_81 :                    
                    7'bzzzzzzz;   
assign sw_output_65 = (control_signal[1] == 0) ? stationary_signal_2:
                      (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :   
                      
                    (control_signal[0] ==0&& index_1 == 7'b1000001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1000001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1000001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1000001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1000001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1000001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1000001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1000001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1000001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1000001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1000001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1000001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1000001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1000001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1000001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1000001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1000001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1000001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1000001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1000001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1000001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1000001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1000001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1000001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1000001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1000001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1000001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1000001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1000001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1000001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1000001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1000001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1000001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1000001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1000001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1000001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1000001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1000001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1000001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1000001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1000001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1000001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1000001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1000001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1000001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1000001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1000001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1000001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1000001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1000001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1000001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1000001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1000001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1000001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1000001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1000001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1000001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1000001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1000001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1000001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1000001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1000001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1000001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1000001) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1000001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1000001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1000001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1000001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1000001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1000001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1000001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1000001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1000001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1000001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1000001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1000001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1000001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1000001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1000001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1000001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000001) ? sw_input_81 :                      
                    7'bzzzzzzz; 
assign sw_output_66 = (control_signal[1] == 0) ? stationary_signal_3:                   
                      (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :  
                      
                    (control_signal[0] ==0&& index_1 == 7'b1000010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1000010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1000010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1000010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1000010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1000010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1000010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1000010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1000010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1000010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1000010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1000010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1000010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1000010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1000010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1000010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1000010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1000010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1000010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1000010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1000010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1000010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1000010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1000010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1000010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1000010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1000010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1000010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1000010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1000010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1000010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1000010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1000010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1000010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1000010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1000010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1000010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1000010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1000010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1000010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1000010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1000010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1000010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1000010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1000010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1000010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1000010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1000010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1000010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1000010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1000010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1000010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1000010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1000010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1000010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1000010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1000010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1000010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1000010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1000010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1000010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1000010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1000010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1000010) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1000010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1000010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1000010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1000010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1000010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1000010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1000010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1000010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1000010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1000010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1000010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1000010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1000010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1000010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1000010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1000010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000010) ? sw_input_81 :                          
                    7'bzzzzzzz; 
assign sw_output_67 = (control_signal[1] == 0) ? stationary_signal_4:
                      (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :   
                      
                    (control_signal[0] ==0&& index_1 == 7'b1000011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1000011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1000011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1000011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1000011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1000011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1000011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1000011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1000011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1000011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1000011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1000011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1000011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1000011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1000011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1000011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1000011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1000011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1000011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1000011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1000011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1000011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1000011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1000011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1000011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1000011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1000011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1000011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1000011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1000011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1000011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1000011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1000011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1000011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1000011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1000011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1000011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1000011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1000011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1000011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1000011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1000011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1000011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1000011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1000011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1000011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1000011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1000011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1000011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1000011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1000011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1000011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1000011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1000011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1000011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1000011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1000011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1000011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1000011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1000011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1000011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1000011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1000011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1000011) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1000011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1000011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1000011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1000011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1000011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1000011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1000011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1000011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1000011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1000011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1000011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1000011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1000011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1000011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1000011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1000011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000011) ? sw_input_81 :           
                    7'bzzzzzzz; 
assign sw_output_68 = (control_signal[1] == 0) ? stationary_signal_5:
                      (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :   
                      
                    (control_signal[0] ==0&& index_1 ==7'b1000100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 ==7'b1000100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 ==7'b1000100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 ==7'b1000100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 ==7'b1000100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 ==7'b1000100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 ==7'b1000100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 ==7'b1000100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 ==7'b1000100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 ==7'b1000100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 ==7'b1000100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 ==7'b1000100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 ==7'b1000100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 ==7'b1000100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 ==7'b1000100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 ==7'b1000100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 ==7'b1000100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 ==7'b1000100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 ==7'b1000100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 ==7'b1000100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 ==7'b1000100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 ==7'b1000100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 ==7'b1000100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 ==7'b1000100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 ==7'b1000100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 ==7'b1000100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 ==7'b1000100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 ==7'b1000100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 ==7'b1000100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 ==7'b1000100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 ==7'b1000100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 ==7'b1000100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 ==7'b1000100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 ==7'b1000100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 ==7'b1000100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 ==7'b1000100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 ==7'b1000100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 ==7'b1000100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 ==7'b1000100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 ==7'b1000100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 ==7'b1000100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 ==7'b1000100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 ==7'b1000100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 ==7'b1000100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 ==7'b1000100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 ==7'b1000100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 ==7'b1000100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 ==7'b1000100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 ==7'b1000100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 ==7'b1000100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 ==7'b1000100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 ==7'b1000100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 ==7'b1000100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 ==7'b1000100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 ==7'b1000100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 ==7'b1000100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 ==7'b1000100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 ==7'b1000100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 ==7'b1000100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 ==7'b1000100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 ==7'b1000100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 ==7'b1000100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 ==7'b1000100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 ==7'b1000100) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 ==7'b1000100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 ==7'b1000100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 ==7'b1000100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 ==7'b1000100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 ==7'b1000100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 ==7'b1000100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 ==7'b1000100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 ==7'b1000100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 ==7'b1000100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 ==7'b1000100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 ==7'b1000100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 ==7'b1000100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 ==7'b1000100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 ==7'b1000100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 ==7'b1000100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 ==7'b1000100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 ==7'b1000100) ? sw_input_81 :                             
                    7'bzzzzzzz;   
assign sw_output_69 = (control_signal[1] == 0) ? stationary_signal_6:
                      (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :   
                      
                    (control_signal[0] ==0&& index_1 ==7'b1000101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 ==7'b1000101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 ==7'b1000101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 ==7'b1000101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 ==7'b1000101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 ==7'b1000101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 ==7'b1000101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 ==7'b1000101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 ==7'b1000101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 ==7'b1000101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 ==7'b1000101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 ==7'b1000101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 ==7'b1000101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 ==7'b1000101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 ==7'b1000101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 ==7'b1000101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 ==7'b1000101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 ==7'b1000101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 ==7'b1000101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 ==7'b1000101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 ==7'b1000101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 ==7'b1000101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 ==7'b1000101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 ==7'b1000101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 ==7'b1000101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 ==7'b1000101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 ==7'b1000101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 ==7'b1000101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 ==7'b1000101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 ==7'b1000101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 ==7'b1000101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 ==7'b1000101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 ==7'b1000101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 ==7'b1000101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 ==7'b1000101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 ==7'b1000101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 ==7'b1000101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 ==7'b1000101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 ==7'b1000101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 ==7'b1000101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 ==7'b1000101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 ==7'b1000101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 ==7'b1000101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 ==7'b1000101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 ==7'b1000101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 ==7'b1000101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 ==7'b1000101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 ==7'b1000101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 ==7'b1000101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 ==7'b1000101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 ==7'b1000101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 ==7'b1000101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 ==7'b1000101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 ==7'b1000101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 ==7'b1000101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 ==7'b1000101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 ==7'b1000101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 ==7'b1000101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 ==7'b1000101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 ==7'b1000101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 ==7'b1000101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 ==7'b1000101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 ==7'b1000101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 ==7'b1000101) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 ==7'b1000101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 ==7'b1000101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 ==7'b1000101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 ==7'b1000101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 ==7'b1000101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 ==7'b1000101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 ==7'b1000101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 ==7'b1000101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 ==7'b1000101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 ==7'b1000101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 ==7'b1000101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 ==7'b1000101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 ==7'b1000101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 ==7'b1000101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 ==7'b1000101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 ==7'b1000101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000101) ? sw_input_81 :                                    
                    7'bzzzzzzz; 
assign sw_output_70 = (control_signal[1] == 0) ? stationary_signal_7:
                      (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :  
                      
                    (control_signal[0] ==0&& index_1 == 7'b1000110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1000110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1000110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1000110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1000110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1000110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1000110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1000110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1000110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1000110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1000110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1000110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1000110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1000110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1000110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1000110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1000110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1000110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1000110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1000110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1000110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1000110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1000110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1000110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1000110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1000110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1000110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1000110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1000110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1000110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1000110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1000110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1000110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1000110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1000110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1000110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1000110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1000110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1000110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1000110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1000110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1000110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1000110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1000110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1000110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1000110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1000110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1000110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1000110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1000110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1000110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1000110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1000110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1000110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1000110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1000110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1000110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1000110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1000110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1000110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1000110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1000110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1000110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1000110) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1000110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1000110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1000110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1000110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1000110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1000110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1000110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1000110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1000110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1000110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1000110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1000110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1000110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1000110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1000110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1000110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000110) ? sw_input_81 :                                  
                    7'bzzzzzzz;    
assign sw_output_71 = (control_signal[1] == 0) ? stationary_signal_8:
                      (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :  
                     
                    (control_signal[0] ==0&& index_1 == 7'b1000111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1000111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1000111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1000111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1000111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1000111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1000111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1000111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1000111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1000111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1000111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1000111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1000111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1000111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1000111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1000111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1000111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1000111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1000111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1000111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1000111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1000111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1000111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1000111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1000111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1000111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1000111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1000111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1000111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1000111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1000111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1000111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1000111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1000111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1000111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1000111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1000111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1000111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1000111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1000111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1000111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1000111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1000111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1000111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1000111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1000111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1000111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1000111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1000111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1000111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1000111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1000111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1000111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1000111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1000111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1000111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1000111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1000111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1000111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1000111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1000111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1000111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1000111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1000111) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1000111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1000111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1000111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1000111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1000111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1000111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1000111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1000111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1000111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1000111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1000111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1000111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1000111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1000111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1000111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1000111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000111) ? sw_input_81 :                       
                    7'bzzzzzzz; 
assign sw_output_72 = (control_signal[1] == 0) ? stationary_signal_9: 
                      (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :   
                      
                    (control_signal[0] ==0&& index_1 == 7'b1001000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001000) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001000) ? sw_input_81 :                          
                    7'bzzzzzzz; 
assign sw_output_73 = (control_signal[1] == 0) ? stationary_signal_1:
                      (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b1001001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001001) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001001) ? sw_input_81 : 
                    7'bzzzzzzz; 
assign sw_output_74 = (control_signal[1] == 0) ? stationary_signal_2:
                      (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :  
                     
                    (control_signal[0] ==0&& index_1 == 7'b1001010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001010) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001010) ? sw_input_81 :                       
                     7'bzzzzzzz;   
assign sw_output_75 = (control_signal[1] == 0) ? stationary_signal_3:
                      (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :  
                      
                    (control_signal[0] ==0&& index_1 == 7'b1001011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001011) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001011) ? sw_input_81 :                     
                     7'bzzzzzzz; 
assign sw_output_76 = (control_signal[1] == 0) ? stationary_signal_4:
                      (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :  
                      
                    (control_signal[0] ==0&& index_1 == 7'b1001100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001100) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001100) ? sw_input_81 :                        
                    7'bzzzzzzz;                         
assign sw_output_77 = (control_signal[1] == 0) ? stationary_signal_5:
                      (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b1001101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001101) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001101) ? sw_input_81 :                       
                    7'bzzzzzzz; 
assign sw_output_78 = (control_signal[1] == 0) ? stationary_signal_6:
                      (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :  
                      
                    (control_signal[0] ==0&& index_1 == 7'b1001110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001110) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001110) ? sw_input_81 :                        
                    7'bzzzzzzz; 
assign sw_output_79 = (control_signal[1] == 0) ? stationary_signal_7:
                      (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 : 
                     
                    (control_signal[0] ==0&& index_1 == 7'b1001111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001111) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001111) ? sw_input_81 : 
                    7'bzzzzzzz; 
assign sw_output_80 = (control_signal[1] == 0) ? stationary_signal_8:
                      (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 : 
                     
                    (control_signal[0] ==0&& index_1 == 7'b1010000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1010000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1010000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1010000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1010000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1010000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1010000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1010000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1010000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1010000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1010000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1010000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1010000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1010000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1010000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1010000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1010000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1010000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1010000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1010000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1010000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1010000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1010000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1010000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1010000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1010000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1010000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1010000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1010000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1010000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1010000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1010000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1010000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1010000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1010000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1010000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1010000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1010000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1010000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1010000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1010000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1010000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1010000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1010000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1010000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1010000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1010000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1010000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1010000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1010000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1010000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1010000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1010000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1010000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1010000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1010000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1010000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1010000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1010000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1010000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1010000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1010000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1010000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1010000) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1010000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1010000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1010000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1010000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1010000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1010000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1010000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1010000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1010000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1010000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1010000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1010000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1010000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1010000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1010000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1010000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1010000) ? sw_input_81 :                     
                    7'bzzzzzzz;   
assign sw_output_81 = (control_signal[1] == 0) ? stationary_signal_9:
                      (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :  
                      
                    (control_signal[0] ==0&& index_1 == 7'b1010001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1010001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1010001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1010001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1010001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1010001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1010001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1010001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1010001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1010001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1010001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1010001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1010001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1010001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1010001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1010001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1010001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1010001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1010001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1010001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1010001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1010001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1010001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1010001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1010001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1010001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1010001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1010001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1010001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1010001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1010001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1010001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1010001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1010001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1010001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1010001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1010001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1010001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1010001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1010001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1010001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1010001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1010001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1010001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1010001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1010001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1010001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1010001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1010001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1010001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1010001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1010001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1010001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1010001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1010001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1010001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1010001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1010001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1010001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1010001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1010001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1010001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1010001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1010001) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1010001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1010001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1010001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1010001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1010001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1010001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1010001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1010001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1010001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1010001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1010001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1010001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1010001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1010001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1010001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1010001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1010001) ? sw_input_81 :                     
                    7'bzzzzzzz; 
assign sw_output_82 = (control_signal[1] == 1) ? stationary_signal_1:
                      (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0000001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0000001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0000001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0000001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0000001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0000001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0000001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0000001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0000001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0000001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0000001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0000001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0000001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0000001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0000001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0000001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0000001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0000001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0000001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0000001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0000001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0000001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0000001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0000001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0000001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0000001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0000001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0000001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0000001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0000001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0000001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0000001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0000001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0000001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0000001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0000001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0000001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0000001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0000001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0000001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0000001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0000001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0000001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0000001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0000001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0000001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0000001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0000001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0000001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0000001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0000001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0000001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0000001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0000001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0000001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0000001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0000001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0000001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0000001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0000001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0000001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0000001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0000001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0000001) ? sw_input_64 :   
                    (control_signal[0] ==0&& index_65 == 7'b0000001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0000001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0000001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0000001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0000001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0000001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0000001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0000001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0000001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0000001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0000001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0000001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0000001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0000001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0000001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0000001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0000001) ? sw_input_81 :                           
                    7'bzzzzzzz;                         
assign sw_output_83 = (control_signal[1] == 1) ? stationary_signal_2:
                      (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 :  
                      
                    (control_signal[0] ==0&& index_1 == 7'b0000010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0000010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0000010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0000010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0000010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0000010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0000010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0000010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0000010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0000010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0000010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0000010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0000010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0000010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0000010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0000010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0000010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0000010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0000010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0000010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0000010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0000010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0000010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0000010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0000010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0000010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0000010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0000010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0000010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0000010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0000010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0000010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0000010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0000010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0000010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0000010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0000010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0000010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0000010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0000010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0000010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0000010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0000010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0000010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0000010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0000010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0000010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0000010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0000010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0000010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0000010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0000010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0000010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0000010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0000010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0000010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0000010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0000010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0000010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0000010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0000010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0000010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0000010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0000010) ? sw_input_64 : 
                     (control_signal[0] ==0&& index_65 == 7'b0000010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0000010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0000010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0000010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0000010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0000010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0000010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0000010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0000010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0000010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0000010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0000010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0000010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0000010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0000010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0000010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0000010) ? sw_input_81 :                        
                    7'bzzzzzzz; 
assign sw_output_84 = (control_signal[1] == 1) ? stationary_signal_3:
                      (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :                     
                      (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0000011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0000011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0000011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0000011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0000011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0000011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0000011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0000011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0000011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0000011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0000011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0000011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0000011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0000011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0000011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0000011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0000011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0000011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0000011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0000011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0000011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0000011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0000011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0000011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0000011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0000011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0000011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0000011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0000011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0000011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0000011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0000011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0000011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0000011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0000011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0000011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0000011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0000011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0000011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0000011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0000011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0000011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0000011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0000011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0000011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0000011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0000011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0000011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0000011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0000011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0000011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0000011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0000011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0000011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0000011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0000011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0000011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0000011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0000011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0000011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0000011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0000011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0000011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0000011) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0000011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0000011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0000011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0000011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0000011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0000011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0000011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0000011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0000011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0000011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0000011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0000011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0000011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0000011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0000011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0000011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0000011) ? sw_input_81 :                       
                     7'bzzzzzzz; 
assign sw_output_85 = (control_signal[1] == 1) ? stationary_signal_4:
                      (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0000100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0000100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0000100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0000100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0000100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0000100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0000100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0000100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0000100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0000100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0000100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0000100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0000100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0000100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0000100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0000100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0000100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0000100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0000100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0000100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0000100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0000100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0000100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0000100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0000100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0000100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0000100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0000100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0000100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0000100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0000100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0000100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0000100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0000100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0000100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0000100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0000100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0000100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0000100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0000100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0000100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0000100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0000100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0000100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0000100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0000100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0000100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0000100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0000100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0000100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0000100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0000100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0000100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0000100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0000100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0000100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0000100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0000100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0000100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0000100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0000100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0000100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0000100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0000100) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0000100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0000100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0000100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0000100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0000100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0000100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0000100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0000100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0000100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0000100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0000100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0000100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0000100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0000100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0000100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0000100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0000100) ? sw_input_81 : 
                     7'bzzzzzzz; 
assign sw_output_86 = (control_signal[1] == 1) ? stationary_signal_5:
                      (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0000101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0000101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0000101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0000101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0000101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0000101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0000101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0000101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0000101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0000101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0000101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0000101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0000101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0000101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0000101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0000101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0000101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0000101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0000101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0000101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0000101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0000101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0000101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0000101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0000101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0000101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0000101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0000101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0000101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0000101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0000101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0000101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0000101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0000101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0000101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0000101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0000101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0000101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0000101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0000101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0000101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0000101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0000101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0000101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0000101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0000101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0000101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0000101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0000101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0000101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0000101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0000101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0000101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0000101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0000101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0000101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0000101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0000101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0000101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0000101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0000101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0000101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0000101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0000101) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0000101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0000101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0000101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0000101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0000101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0000101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0000101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0000101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0000101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0000101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0000101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0000101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0000101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0000101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0000101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0000101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0000101) ? sw_input_81 :                   
                    7'bzzzzzzz;   
assign sw_output_87 = (control_signal[1] == 1) ? stationary_signal_6:
                      (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0000110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0000110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0000110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0000110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0000110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0000110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0000110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0000110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0000110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0000110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0000110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0000110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0000110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0000110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0000110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0000110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0000110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0000110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0000110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0000110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0000110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0000110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0000110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0000110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0000110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0000110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0000110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0000110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0000110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0000110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0000110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0000110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0000110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0000110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0000110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0000110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0000110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0000110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0000110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0000110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0000110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0000110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0000110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0000110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0000110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0000110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0000110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0000110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0000110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0000110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0000110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0000110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0000110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0000110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0000110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0000110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0000110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0000110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0000110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0000110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0000110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0000110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0000110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0000110) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0000110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0000110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0000110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0000110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0000110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0000110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0000110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0000110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0000110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0000110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0000110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0000110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0000110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0000110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0000110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0000110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0000110) ? sw_input_81 :                       
                     7'bzzzzzzz; 
assign sw_output_88 = (control_signal[1] == 1) ? stationary_signal_7:
                      (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 :  
                      
                    (control_signal[0] ==0&& index_1 == 7'b0000111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0000111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0000111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0000111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0000111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0000111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0000111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0000111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0000111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0000111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0000111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0000111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0000111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0000111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0000111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0000111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0000111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0000111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0000111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0000111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0000111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0000111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0000111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0000111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0000111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0000111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0000111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0000111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0000111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0000111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0000111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0000111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0000111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0000111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0000111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0000111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0000111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0000111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0000111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0000111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0000111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0000111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0000111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0000111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0000111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0000111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0000111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0000111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0000111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0000111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0000111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0000111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0000111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0000111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0000111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0000111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0000111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0000111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0000111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0000111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0000111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0000111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0000111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0000111) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0000111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0000111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0000111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0000111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0000111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0000111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0000111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0000111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0000111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0000111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0000111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0000111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0000111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0000111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0000111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0000111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0000111) ? sw_input_81 :                                                                  
                     7'bzzzzzzz;                         
assign sw_output_89 = (control_signal[1] == 1) ? stationary_signal_8:
                      (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :                     
                      (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001000) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0001000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001000) ? sw_input_81 :                         
                     7'bzzzzzzz; 
assign sw_output_90 = (control_signal[1] == 1) ? stationary_signal_9:
                      (control_signal[0] ==1&& index_1 == 7'b0000001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000001) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000001) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000001) ? sw_input_9 :  
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001001) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0001001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001001) ? sw_input_81 :                     
                    7'bzzzzzzz; 
assign sw_output_91 = (control_signal[1] == 1) ? stationary_signal_10:
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001010) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0001010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001010) ? sw_input_81 :  
                    7'bzzzzzzz; 
assign sw_output_92 = (control_signal[1] == 1) ? stationary_signal_11:
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001011) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0001011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001011) ? sw_input_81 :                   
                     7'bzzzzzzz;   
assign sw_output_93 = (control_signal[1] == 1) ? stationary_signal_12:
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :                     
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001100) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0001100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001100) ? sw_input_81 :                       
                    7'bzzzzzzz; 
assign sw_output_94 = (control_signal[1] == 1) ? stationary_signal_13:
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :                     
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001101) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0001101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001101) ? sw_input_81 :                                              
                    7'bzzzzzzz;                         
assign sw_output_95 = (control_signal[1] == 1) ? stationary_signal_14: 
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001110) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0001110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001110) ? sw_input_81 :                        
                     7'bzzzzzzz; 
assign sw_output_96 = (control_signal[1] == 1) ? stationary_signal_15:
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0001111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0001111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0001111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0001111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0001111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0001111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0001111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0001111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0001111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0001111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0001111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0001111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0001111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0001111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0001111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0001111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0001111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0001111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0001111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0001111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0001111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0001111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0001111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0001111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0001111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0001111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0001111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0001111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0001111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0001111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0001111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0001111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0001111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0001111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0001111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0001111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0001111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0001111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0001111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0001111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0001111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0001111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0001111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0001111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0001111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0001111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0001111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0001111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0001111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0001111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0001111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0001111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0001111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0001111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0001111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0001111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0001111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0001111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0001111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0001111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0001111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0001111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0001111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0001111) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0001111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0001111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0001111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0001111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0001111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0001111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0001111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0001111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0001111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0001111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0001111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0001111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0001111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0001111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0001111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0001111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0001111) ? sw_input_81 :                          
                    7'bzzzzzzz; 
assign sw_output_97 = (control_signal[1] == 1) ? stationary_signal_16:
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0010000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010000) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0010000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010000) ? sw_input_81 : 
                    7'bzzzzzzz; 
assign sw_output_98 = (control_signal[1] == 1) ? stationary_signal_17:
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 :  
                      
                    (control_signal[0] ==0&& index_1 == 7'b0010001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010001) ? sw_input_64 :
                     (control_signal[0] ==0&& index_65 == 7'b0010001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010001) ? sw_input_81 :                     
                     7'bzzzzzzz;   
assign sw_output_99 = (control_signal[1] == 1) ? stationary_signal_18:
                      (control_signal[0] ==1&& index_1 == 7'b0000010) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000010) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000010) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000010) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000010) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000010) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000010) ? sw_input_7 :
                      (control_signal[0] ==1&& index_8 == 7'b0000010) ? sw_input_8 :                      
                      (control_signal[0] ==1&& index_9 == 7'b0000010) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0010010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010010) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0010010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010010) ? sw_input_81 :                       
                    7'bzzzzzzz; 
assign sw_output_100 =(control_signal[1] == 1) ? stationary_signal_19:
                      (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0010011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010011) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0010011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010011) ? sw_input_81 :                          
                    7'bzzzzzzz;                         
assign sw_output_101 =(control_signal[1] == 1) ? stationary_signal_20:
                      (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 : 
                      
                    (control_signal[0] ==0&& index_1 == 7'b0010100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010100) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0010100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010100) ? sw_input_81 :                       
                    7'bzzzzzzz; 
assign sw_output_102 =(control_signal[1] == 1) ? stationary_signal_21:
                     
                          (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 : 
                      
                       (control_signal[0] ==0&& index_1 == 7'b0010101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010101) ? sw_input_64 :
                     (control_signal[0] ==0&& index_65 == 7'b0010101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010101) ? sw_input_81 :                        
                      7'bzzzzzzz; 
assign sw_output_103 =(control_signal[1] == 1) ? stationary_signal_22:
                      
                       (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 :
                      
                       (control_signal[0] ==0&& index_1 == 7'b0010110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010110) ? sw_input_64 : 
                     (control_signal[0] ==0&& index_65 == 7'b0010110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010110) ? sw_input_81 :
                      7'bzzzzzzz; 
assign sw_output_104 =(control_signal[1] == 1) ? stationary_signal_23:
                     
                         (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 : 
                     
                       (control_signal[0] ==0&& index_1 == 7'b0010111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0010111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0010111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0010111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0010111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0010111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0010111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0010111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0010111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0010111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0010111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0010111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0010111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0010111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0010111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0010111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0010111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0010111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0010111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0010111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0010111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0010111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0010111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0010111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0010111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0010111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0010111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0010111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0010111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0010111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0010111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0010111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0010111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0010111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0010111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0010111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0010111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0010111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0010111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0010111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0010111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0010111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0010111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0010111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0010111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0010111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0010111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0010111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0010111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0010111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0010111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0010111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0010111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0010111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0010111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0010111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0010111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0010111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0010111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0010111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0010111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0010111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0010111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0010111) ? sw_input_64 :
                     (control_signal[0] ==0&& index_65 == 7'b0010111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0010111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0010111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0010111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0010111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0010111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0010111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0010111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0010111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0010111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0010111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0010111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0010111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0010111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0010111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0010111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0010111) ? sw_input_81 :                   
                      7'bzzzzzzz;   
assign sw_output_105 = (control_signal[1] == 1) ? stationary_signal_24:
                     
                         (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 : 
                      
                      (control_signal[0] ==0&& index_1 == 7'b0011000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011000) ? sw_input_64 : 
                     (control_signal[0] ==0&& index_65 == 7'b0011000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011000) ? sw_input_81 :                       
                      7'bzzzzzzz; 
assign sw_output_106 =(control_signal[1] == 1) ? stationary_signal_25:
                      
                        (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 :
                      
                     (control_signal[0] ==0&& index_1 == 7'b0011001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011001) ? sw_input_64 : 
                     (control_signal[0] ==0&& index_65 == 7'b0011001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011001) ? sw_input_81 :                       
                      7'bzzzzzzz;                         
assign sw_output_107 =(control_signal[1] == 1) ? stationary_signal_26:
                     
                         (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 : 
                       
                       (control_signal[0] ==0&& index_1 == 7'b0011010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011010) ? sw_input_64 :
                     (control_signal[0] ==0&& index_65 == 7'b0011010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011010) ? sw_input_81 :                       
                     7'bzzzzzzz; 
assign sw_output_108 = (control_signal[1] == 1) ? stationary_signal_27:
                      
                         (control_signal[0] ==1&& index_1 == 7'b0000011) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000011) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000011) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000011) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000011) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000011) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000011) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000011) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000011) ? sw_input_9 :
                      
                      (control_signal[0] ==0&& index_1 == 7'b0011011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011011) ? sw_input_64 :
                     (control_signal[0] ==0&& index_65 == 7'b0011011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011011) ? sw_input_81 :                      
                      7'bzzzzzzz; 
assign sw_output_109 =(control_signal[1] == 1) ? stationary_signal_28:
                     
                      (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :
                      
                      (control_signal[0] ==0&& index_1 == 7'b0011100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011100) ? sw_input_64 :
                     (control_signal[0] ==0&& index_65 == 7'b0011100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011100) ? sw_input_81 : 
                      7'bzzzzzzz; 
assign sw_output_110 =(control_signal[1] == 1) ? stationary_signal_29:
                     
                        (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 : 
                      
                      (control_signal[0] ==0&& index_1 == 7'b0011101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011101) ? sw_input_64 :
                     (control_signal[0] ==0&& index_65 == 7'b0011101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011101) ? sw_input_81 :                    
                      7'bzzzzzzz;   
assign sw_output_111 =(control_signal[1] == 1) ? stationary_signal_30:
                      
                        (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :
                     
                      (control_signal[0] ==0&& index_1 == 7'b0011110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011110) ? sw_input_64 :
                     (control_signal[0] ==0&& index_65 == 7'b0011110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011110) ? sw_input_81 :                      
                      7'bzzzzzzz; 
assign sw_output_112 =(control_signal[1] == 1) ? stationary_signal_31:
                     
                        (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 : 
                      
                      (control_signal[0] ==0&& index_1 == 7'b0011111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0011111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0011111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0011111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0011111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0011111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0011111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0011111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0011111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0011111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0011111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0011111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0011111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0011111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0011111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0011111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0011111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0011111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0011111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0011111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0011111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0011111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0011111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0011111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0011111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0011111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0011111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0011111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0011111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0011111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0011111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0011111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0011111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0011111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0011111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0011111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0011111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0011111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0011111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0011111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0011111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0011111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0011111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0011111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0011111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0011111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0011111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0011111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0011111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0011111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0011111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0011111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0011111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0011111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0011111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0011111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0011111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0011111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0011111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0011111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0011111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0011111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0011111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0011111) ? sw_input_64 :
                     (control_signal[0] ==0&& index_65 == 7'b0011111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0011111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0011111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0011111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0011111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0011111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0011111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0011111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0011111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0011111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0011111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0011111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0011111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0011111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0011111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0011111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0011111) ? sw_input_81 :                      
                      7'bzzzzzzz;                         
assign sw_output_113 =(control_signal[1] == 1) ? stationary_signal_32: 
                  
                        (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 : 
                      
                      (control_signal[0] ==0&& index_1 == 7'b0100000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100000) ? sw_input_64 : 
                     (control_signal[0] ==0&& index_65 == 7'b0100000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100000) ? sw_input_81 :                       
                     7'bzzzzzzz; 
assign sw_output_114 = (control_signal[1] == 1) ? stationary_signal_33:
                     
                         (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :  
                      
                       (control_signal[0] ==0&& index_1 == 7'b0100001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100001) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100001) ? sw_input_81 :                   
                      7'bzzzzzzz; 
assign sw_output_115 =(control_signal[1] == 1) ? stationary_signal_34:
                     
                         (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 : 
                      
                        (control_signal[0] ==0&& index_1 == 7'b0100010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100010) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100010) ? sw_input_81 :
                      7'bzzzzzzz; 
assign sw_output_116 =(control_signal[1] == 1) ? stationary_signal_35:
                     
                         (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :
                      
                     (control_signal[0] ==0&& index_1 == 7'b0100011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100011) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100011) ? sw_input_81 :
                                       
                      7'bzzzzzzz;   
assign sw_output_117 =(control_signal[1] == 1) ? stationary_signal_36:
                     
                        (control_signal[0] ==1&& index_1 == 7'b0000100) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000100) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000100) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000100) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000100) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000100) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000100) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000100) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000100) ? sw_input_9 :
                      
                      (control_signal[0] ==0&& index_1 == 7'b0100100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100100) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100100) ? sw_input_81 :                      
                      7'bzzzzzzz; 
assign sw_output_118 =(control_signal[1] == 1) ? stationary_signal_37:
                     
                        (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 : 
                      
         
                      
                       (control_signal[0] ==0&& index_1 == 7'b0100101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100101) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100101) ? sw_input_81 :                      
                      7'bzzzzzzz;                         
assign sw_output_119 =(control_signal[1] == 1) ? stationary_signal_38:
                     
                         (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 : 
                      
                        (control_signal[0] ==0&& index_1 == 7'b0100110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100110) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100110) ? sw_input_81 :                      
                     7'bzzzzzzz; 
assign sw_output_120 =(control_signal[1] == 1) ? stationary_signal_39:                   
                       
                         (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 : 
                      
                        (control_signal[0] ==0&& index_1 == 7'b0100111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0100111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0100111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0100111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0100111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0100111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0100111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0100111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0100111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0100111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0100111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0100111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0100111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0100111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0100111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0100111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0100111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0100111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0100111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0100111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0100111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0100111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0100111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0100111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0100111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0100111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0100111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0100111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0100111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0100111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0100111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0100111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0100111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0100111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0100111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0100111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0100111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0100111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0100111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0100111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0100111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0100111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0100111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0100111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0100111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0100111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0100111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0100111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0100111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0100111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0100111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0100111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0100111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0100111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0100111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0100111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0100111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0100111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0100111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0100111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0100111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0100111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0100111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0100111) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0100111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0100111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0100111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0100111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0100111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0100111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0100111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0100111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0100111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0100111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0100111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0100111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0100111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0100111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0100111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0100111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0100111) ? sw_input_81 :                        
                      7'bzzzzzzz; 
assign sw_output_121 =(control_signal[1] == 1) ? stationary_signal_40:                   
                        (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 : 
                      
                        (control_signal[0] ==0&& index_1 == 7'b0101000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101000) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101000) ? sw_input_81 : 
                      7'bzzzzzzz; 
assign sw_output_122 =(control_signal[1] == 1) ? stationary_signal_41:                 
                       (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 :
                     
                      (control_signal[0] ==0&& index_1 == 7'b0101001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101001) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101001) ? sw_input_81 :                      
                      7'bzzzzzzz;   
assign sw_output_123 =(control_signal[1] == 1) ? stationary_signal_42:             
                       (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 : 
                      
                      (control_signal[0] ==0&& index_1 == 7'b0101010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101010) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101010) ? sw_input_81 :                        
                      7'bzzzzzzz; 
assign sw_output_124 =(control_signal[1] == 1) ? stationary_signal_43:                    
                          (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 : 
                      
                     (control_signal[0] ==0&& index_1 == 7'b0101011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101011) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101011) ? sw_input_81 :                         
                      7'bzzzzzzz;                         
assign sw_output_125 =(control_signal[1] == 1) ? stationary_signal_44:                    
                         (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 : 
                      
                      (control_signal[0] ==0&& index_1 == 7'b0101100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101100) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101100) ? sw_input_81 :                        
                     7'bzzzzzzz; 
assign sw_output_126 =(control_signal[1] == 1) ? stationary_signal_45:                    
                         (control_signal[0] ==1&& index_1 == 7'b0000101) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000101) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000101) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000101) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000101) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000101) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000101) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000101) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000101) ? sw_input_9 :
                     
                     (control_signal[0] ==0&& index_1 == 7'b0101101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101101) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101101) ? sw_input_81 :                         
                      7'bzzzzzzz; 
assign sw_output_127 =(control_signal[1] == 1) ? stationary_signal_46:                    
                     
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                      
                       (control_signal[0] ==0&& index_1 == 7'b0101110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101110) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101110) ? sw_input_81 : 
                      7'bzzzzzzz; 
assign sw_output_128 =(control_signal[1] == 1) ? stationary_signal_47:   
                
                        (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                      
                      
                     (control_signal[0] ==0&& index_1 == 7'b0101111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0101111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0101111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0101111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0101111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0101111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0101111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0101111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0101111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0101111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0101111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0101111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0101111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0101111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0101111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0101111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0101111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0101111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0101111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0101111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0101111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0101111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0101111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0101111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0101111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0101111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0101111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0101111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0101111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0101111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0101111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0101111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0101111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0101111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0101111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0101111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0101111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0101111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0101111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0101111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0101111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0101111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0101111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0101111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0101111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0101111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0101111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0101111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0101111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0101111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0101111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0101111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0101111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0101111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0101111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0101111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0101111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0101111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0101111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0101111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0101111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0101111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0101111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0101111) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0101111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0101111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0101111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0101111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0101111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0101111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0101111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0101111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0101111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0101111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0101111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0101111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0101111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0101111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0101111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0101111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0101111) ? sw_input_81 :                       
                      7'bzzzzzzz;   
assign sw_output_129 =(control_signal[1] == 1) ? stationary_signal_48:

                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                      
                      
                       
                    
                    (control_signal[0] ==0&& index_1 == 7'b0110000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110000) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110000) ? sw_input_81 :            
                    7'bzzzzzzz; 
 assign sw_output_130 =(control_signal[1] == 1) ? stationary_signal_49:
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                    
                   (control_signal[0] ==0&& index_1 == 7'b0110001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110001) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110001) ? sw_input_81 :           
                    7'bzzzzzzz; 
 assign sw_output_131 =(control_signal[1] == 1) ? stationary_signal_50:
                     (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b0110010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110010) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110010) ? sw_input_81 :            
                    7'bzzzzzzz; 
  assign sw_output_132 =(control_signal[1] == 1) ? stationary_signal_51:
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                    
                     (control_signal[0] ==0&& index_1 == 7'b0110011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110011) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110001) ? sw_input_81 :            
                    7'bzzzzzzz; 
  assign sw_output_133 =(control_signal[1] == 1) ? stationary_signal_52:
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                    
                   (control_signal[0] ==0&& index_1 == 7'b0110100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110100) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110100) ? sw_input_81 :            
                    7'bzzzzzzz; 
assign sw_output_134 =(control_signal[1] == 1) ? stationary_signal_53:
                     (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                    
                    
                    (control_signal[0] ==0&& index_1 == 7'b0110101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110101) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110101) ? sw_input_81 :            
                    7'bzzzzzzz; 
assign sw_output_135 =(control_signal[1] == 1) ? stationary_signal_54:
                      (control_signal[0] ==1&& index_1 == 7'b0000110) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000110) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000110) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000110) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000110) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000110) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000110) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000110) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000110) ? sw_input_9 :
                    
                   (control_signal[0] ==0&& index_1 == 7'b0110110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110110) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110110) ? sw_input_81 :            
                    7'bzzzzzzz; 
assign sw_output_136 =(control_signal[1] == 1) ? stationary_signal_55:
                     (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b0110111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0110111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0110111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0110111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0110111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0110111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0110111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0110111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0110111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0110111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0110111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0110111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0110111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0110111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0110111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0110111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0110111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0110111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0110111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0110111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0110111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0110111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0110111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0110111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0110111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0110111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0110111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0110111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0110111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0110111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0110111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0110111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0110111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0110111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0110111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0110111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0110111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0110111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0110111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0110111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0110111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0110111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0110111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0110111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0110111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0110111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0110111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0110111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0110111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0110111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0110111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0110111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0110111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0110111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0110111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0110111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0110111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0110111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0110111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0110111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0110111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0110111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0110111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0110111) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0110111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0110111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0110111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0110111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0110111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0110111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0110111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0110111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0110111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0110111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0110111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0110111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0110111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0110111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0110111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0110111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0110111) ? sw_input_81 :            
                    7'bzzzzzzz; 
  assign sw_output_137 =(control_signal[1] == 1) ? stationary_signal_56:
                     (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b0111000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111000) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0111000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111000) ? sw_input_81 :            
                    7'bzzzzzzz; 
assign sw_output_138 =(control_signal[1] == 1) ? stationary_signal_57:
                     (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                    
                   (control_signal[0] ==0&& index_1 == 7'b0111001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111001) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0111001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111001) ? sw_input_81 :            
                    7'bzzzzzzz; 
  assign sw_output_139 =(control_signal[1] == 1) ? stationary_signal_58:
                     (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b0111010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111010) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0111010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111010) ? sw_input_81 :           
                    7'bzzzzzzz; 
  assign sw_output_140 =(control_signal[1] == 1) ? stationary_signal_59:
                    (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b0111011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111011) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0111011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111011) ? sw_input_81 :             
                    7'bzzzzzzz; 
assign sw_output_141 =(control_signal[1] == 1) ? stationary_signal_60:
                     (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                    
                   (control_signal[0] ==0&& index_1 == 7'b0111100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111100) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0111100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111100) ? sw_input_81 :            
                    7'bzzzzzzz; 
 assign sw_output_142 =(control_signal[1] == 1) ? stationary_signal_61:
                    (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                    
                     (control_signal[0] ==0&& index_1 == 7'b0111101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111101) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0111101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111101) ? sw_input_81 :            
                    7'bzzzzzzz; 
assign sw_output_143 =(control_signal[1] == 1) ? stationary_signal_62:
                    (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b0111110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111110) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b0111110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111110) ? sw_input_81 : 
                    
                                  
                    7'bzzzzzzz; 
assign sw_output_144 =(control_signal[1] == 1) ? stationary_signal_63:
                      (control_signal[0] ==1&& index_1 == 7'b0000111) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0000111) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0000111) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0000111) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0000111) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0000111) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0000111) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0000111) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0000111) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b0111111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b0111111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b0111111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b0111111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b0111111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b0111111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b0111111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b0111111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b0111111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b0111111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b0111111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b0111111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b0111111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b0111111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b0111111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b0111111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b0111111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b0111111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b0111111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b0111111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b0111111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b0111111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b0111111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b0111111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b0111111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b0111111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b0111111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b0111111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b0111111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b0111111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b0111111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b0111111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b0111111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b0111111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b0111111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b0111111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b0111111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b0111111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b0111111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b0111111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b0111111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b0111111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b0111111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b0111111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b0111111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b0111111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b0111111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b0111111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b0111111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b0111111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b0111111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b0111111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b0111111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b0111111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b0111111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b0111111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b0111111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b0111111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b0111111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b0111111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b0111111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b0111111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b0111111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b0111111) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b0111111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b0111111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b0111111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b0111111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b0111111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b0111111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b0111111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b0111111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b0111111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b0111111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b0111111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b0111111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b0111111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b0111111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b0111111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b0111111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b0111111) ? sw_input_81 :           
                    7'bzzzzzzz; 
assign sw_output_145 =(control_signal[1] == 1) ? stationary_signal_64:
                    (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b1000000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1000000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1000000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1000000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1000000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1000000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1000000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1000000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1000000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1000000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1000000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1000000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1000000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1000000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1000000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1000000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1000000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1000000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1000000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1000000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1000000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1000000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1000000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1000000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1000000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1000000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1000000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1000000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1000000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1000000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1000000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1000000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1000000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1000000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1000000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1000000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1000000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1000000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1000000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1000000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1000000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1000000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1000000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1000000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1000000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1000000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1000000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1000000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1000000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1000000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1000000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1000000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1000000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1000000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1000000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1000000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1000000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1000000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1000000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1000000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1000000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1000000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1000000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1000000) ? sw_input_64 :
                    (control_signal[0] ==0&& index_65 == 7'b1000000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1000000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1000000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1000000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1000000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1000000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1000000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1000000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1000000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1000000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1000000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1000000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1000000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1000000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1000000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1000000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000000) ? sw_input_81 :            
                    7'bzzzzzzz; 
assign sw_output_146 =(control_signal[1] == 1) ? stationary_signal_65:

                    (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :
                      
                    (control_signal[0] ==0&& index_1 == 7'b1000001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1000001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1000001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1000001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1000001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1000001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1000001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1000001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1000001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1000001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1000001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1000001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1000001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1000001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1000001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1000001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1000001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1000001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1000001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1000001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1000001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1000001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1000001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1000001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1000001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1000001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1000001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1000001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1000001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1000001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1000001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1000001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1000001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1000001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1000001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1000001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1000001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1000001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1000001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1000001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1000001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1000001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1000001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1000001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1000001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1000001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1000001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1000001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1000001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1000001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1000001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1000001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1000001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1000001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1000001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1000001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1000001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1000001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1000001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1000001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1000001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1000001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1000001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1000001) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1000001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1000001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1000001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1000001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1000001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1000001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1000001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1000001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1000001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1000001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1000001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1000001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1000001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1000001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1000001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1000001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000001) ? sw_input_81 :            
                    7'bzzzzzzz; 
assign sw_output_147 =(control_signal[1] == 1) ? stationary_signal_66:
                    (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :
                    
                     (control_signal[0] ==0&& index_1 == 7'b1000010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1000010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1000010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1000010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1000010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1000010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1000010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1000010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1000010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1000010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1000010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1000010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1000010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1000010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1000010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1000010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1000010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1000010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1000010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1000010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1000010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1000010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1000010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1000010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1000010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1000010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1000010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1000010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1000010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1000010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1000010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1000010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1000010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1000010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1000010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1000010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1000010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1000010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1000010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1000010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1000010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1000010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1000010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1000010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1000010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1000010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1000010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1000010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1000010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1000010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1000010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1000010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1000010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1000010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1000010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1000010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1000010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1000010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1000010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1000010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1000010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1000010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1000010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1000010) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1000010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1000010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1000010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1000010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1000010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1000010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1000010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1000010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1000010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1000010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1000010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1000010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1000010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1000010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1000010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1000010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000010) ? sw_input_81 :            
                    7'bzzzzzzz; 
  assign sw_output_148 =(control_signal[1] == 1) ? stationary_signal_67:
                    (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b1000011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1000011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1000011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1000011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1000011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1000011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1000011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1000011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1000011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1000011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1000011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1000011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1000011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1000011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1000011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1000011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1000011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1000011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1000011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1000011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1000011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1000011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1000011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1000011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1000011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1000011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1000011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1000011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1000011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1000011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1000011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1000011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1000011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1000011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1000011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1000011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1000011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1000011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1000011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1000011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1000011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1000011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1000011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1000011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1000011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1000011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1000011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1000011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1000011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1000011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1000011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1000011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1000011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1000011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1000011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1000011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1000011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1000011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1000011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1000011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1000011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1000011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1000011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1000011) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1000011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1000011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1000011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1000011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1000011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1000011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1000011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1000011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1000011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1000011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1000011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1000011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1000011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1000011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1000011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1000011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000011) ? sw_input_81 :            
                    7'bzzzzzzz; 
  assign sw_output_149 =(control_signal[1] == 1) ? stationary_signal_68:
                    (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 ==7'b1000100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 ==7'b1000100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 ==7'b1000100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 ==7'b1000100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 ==7'b1000100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 ==7'b1000100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 ==7'b1000100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 ==7'b1000100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 ==7'b1000100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 ==7'b1000100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 ==7'b1000100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 ==7'b1000100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 ==7'b1000100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 ==7'b1000100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 ==7'b1000100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 ==7'b1000100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 ==7'b1000100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 ==7'b1000100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 ==7'b1000100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 ==7'b1000100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 ==7'b1000100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 ==7'b1000100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 ==7'b1000100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 ==7'b1000100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 ==7'b1000100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 ==7'b1000100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 ==7'b1000100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 ==7'b1000100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 ==7'b1000100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 ==7'b1000100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 ==7'b1000100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 ==7'b1000100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 ==7'b1000100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 ==7'b1000100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 ==7'b1000100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 ==7'b1000100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 ==7'b1000100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 ==7'b1000100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 ==7'b1000100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 ==7'b1000100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 ==7'b1000100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 ==7'b1000100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 ==7'b1000100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 ==7'b1000100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 ==7'b1000100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 ==7'b1000100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 ==7'b1000100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 ==7'b1000100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 ==7'b1000100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 ==7'b1000100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 ==7'b1000100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 ==7'b1000100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 ==7'b1000100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 ==7'b1000100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 ==7'b1000100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 ==7'b1000100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 ==7'b1000100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 ==7'b1000100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 ==7'b1000100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 ==7'b1000100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 ==7'b1000100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 ==7'b1000100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 ==7'b1000100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 ==7'b1000100) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 ==7'b1000100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 ==7'b1000100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 ==7'b1000100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 ==7'b1000100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 ==7'b1000100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 ==7'b1000100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 ==7'b1000100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 ==7'b1000100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 ==7'b1000100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 ==7'b1000100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 ==7'b1000100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 ==7'b1000100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 ==7'b1000100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 ==7'b1000100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 ==7'b1000100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 ==7'b1000100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 ==7'b1000100) ? sw_input_81 :            
                    7'bzzzzzzz; 
assign sw_output_150 =(control_signal[1] == 1) ? stationary_signal_69:
                    (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :
                    
                     (control_signal[0] ==0&& index_1 ==7'b1000101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 ==7'b1000101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 ==7'b1000101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 ==7'b1000101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 ==7'b1000101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 ==7'b1000101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 ==7'b1000101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 ==7'b1000101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 ==7'b1000101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 ==7'b1000101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 ==7'b1000101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 ==7'b1000101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 ==7'b1000101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 ==7'b1000101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 ==7'b1000101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 ==7'b1000101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 ==7'b1000101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 ==7'b1000101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 ==7'b1000101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 ==7'b1000101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 ==7'b1000101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 ==7'b1000101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 ==7'b1000101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 ==7'b1000101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 ==7'b1000101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 ==7'b1000101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 ==7'b1000101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 ==7'b1000101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 ==7'b1000101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 ==7'b1000101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 ==7'b1000101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 ==7'b1000101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 ==7'b1000101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 ==7'b1000101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 ==7'b1000101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 ==7'b1000101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 ==7'b1000101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 ==7'b1000101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 ==7'b1000101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 ==7'b1000101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 ==7'b1000101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 ==7'b1000101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 ==7'b1000101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 ==7'b1000101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 ==7'b1000101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 ==7'b1000101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 ==7'b1000101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 ==7'b1000101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 ==7'b1000101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 ==7'b1000101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 ==7'b1000101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 ==7'b1000101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 ==7'b1000101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 ==7'b1000101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 ==7'b1000101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 ==7'b1000101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 ==7'b1000101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 ==7'b1000101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 ==7'b1000101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 ==7'b1000101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 ==7'b1000101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 ==7'b1000101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 ==7'b1000101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 ==7'b1000101) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 ==7'b1000101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 ==7'b1000101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 ==7'b1000101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 ==7'b1000101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 ==7'b1000101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 ==7'b1000101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 ==7'b1000101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 ==7'b1000101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 ==7'b1000101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 ==7'b1000101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 ==7'b1000101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 ==7'b1000101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 ==7'b1000101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 ==7'b1000101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 ==7'b1000101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 ==7'b1000101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000101) ? sw_input_81 :             
                    7'bzzzzzzz; 
assign sw_output_151 =(control_signal[1] == 1) ? stationary_signal_70:
                    (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :
                    
                     (control_signal[0] ==0&& index_1 == 7'b1000110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1000110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1000110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1000110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1000110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1000110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1000110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1000110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1000110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1000110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1000110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1000110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1000110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1000110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1000110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1000110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1000110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1000110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1000110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1000110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1000110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1000110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1000110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1000110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1000110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1000110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1000110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1000110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1000110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1000110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1000110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1000110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1000110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1000110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1000110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1000110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1000110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1000110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1000110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1000110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1000110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1000110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1000110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1000110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1000110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1000110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1000110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1000110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1000110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1000110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1000110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1000110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1000110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1000110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1000110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1000110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1000110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1000110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1000110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1000110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1000110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1000110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1000110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1000110) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1000110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1000110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1000110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1000110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1000110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1000110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1000110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1000110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1000110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1000110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1000110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1000110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1000110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1000110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1000110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1000110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000110) ? sw_input_81 :            
                    7'bzzzzzzz; 
assign sw_output_152 =(control_signal[1] == 1) ? stationary_signal_71:
                    (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :
                    
                     (control_signal[0] ==0&& index_1 == 7'b1000111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1000111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1000111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1000111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1000111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1000111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1000111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1000111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1000111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1000111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1000111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1000111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1000111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1000111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1000111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1000111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1000111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1000111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1000111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1000111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1000111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1000111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1000111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1000111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1000111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1000111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1000111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1000111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1000111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1000111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1000111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1000111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1000111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1000111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1000111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1000111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1000111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1000111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1000111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1000111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1000111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1000111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1000111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1000111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1000111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1000111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1000111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1000111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1000111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1000111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1000111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1000111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1000111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1000111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1000111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1000111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1000111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1000111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1000111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1000111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1000111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1000111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1000111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1000111) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1000111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1000111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1000111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1000111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1000111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1000111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1000111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1000111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1000111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1000111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1000111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1000111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1000111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1000111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1000111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1000111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1000111) ? sw_input_81 :            
                    7'bzzzzzzz; 
 assign sw_output_153 =(control_signal[1] == 1) ? stationary_signal_72:
                      (control_signal[0] ==1&& index_1 == 7'b0001000) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001000) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001000) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001000) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001000) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001000) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001000) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001000) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001000) ? sw_input_9 :
                    
                     (control_signal[0] ==0&& index_1 == 7'b1001000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001000) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001000) ? sw_input_81 :            
                    7'bzzzzzzz; 
assign sw_output_154 =(control_signal[1] == 1) ? stationary_signal_73:
                    (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :
                    
                     (control_signal[0] ==0&& index_1 == 7'b1001001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001001) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001001) ? sw_input_81 :             
                    7'bzzzzzzz; 
   assign sw_output_155 =(control_signal[1] == 1) ? stationary_signal_74:
   
                    (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b1001010) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001010) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001010) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001010) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001010) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001010) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001010) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001010) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001010) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001010) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001010) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001010) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001010) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001010) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001010) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001010) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001010) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001010) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001010) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001010) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001010) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001010) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001010) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001010) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001010) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001010) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001010) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001010) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001010) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001010) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001010) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001010) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001010) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001010) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001010) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001010) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001010) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001010) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001010) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001010) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001010) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001010) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001010) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001010) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001010) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001010) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001010) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001010) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001010) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001010) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001010) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001010) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001010) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001010) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001010) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001010) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001010) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001010) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001010) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001010) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001010) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001010) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001010) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001010) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001010) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001010) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001010) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001010) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001010) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001010) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001010) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001010) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001010) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001010) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001010) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001010) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001010) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001010) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001010) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001010) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001010) ? sw_input_81 :            
                    7'bzzzzzzz; 
  assign sw_output_156 =(control_signal[1] == 1) ? stationary_signal_75:
  
                     (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :
                    
                     (control_signal[0] ==0&& index_1 == 7'b1001011) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001011) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001011) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001011) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001011) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001011) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001011) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001011) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001011) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001011) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001011) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001011) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001011) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001011) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001011) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001011) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001011) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001011) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001011) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001011) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001011) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001011) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001011) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001011) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001011) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001011) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001011) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001011) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001011) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001011) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001011) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001011) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001011) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001011) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001011) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001011) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001011) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001011) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001011) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001011) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001011) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001011) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001011) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001011) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001011) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001011) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001011) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001011) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001011) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001011) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001011) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001011) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001011) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001011) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001011) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001011) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001011) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001011) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001011) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001011) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001011) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001011) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001011) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001011) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001011) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001011) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001011) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001011) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001011) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001011) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001011) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001011) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001011) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001011) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001011) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001011) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001011) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001011) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001011) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001011) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001011) ? sw_input_81 :           
                    7'bzzzzzzz; 
  assign sw_output_157 =(control_signal[1] == 1) ? stationary_signal_76:
  
                     (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b1001100) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001100) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001100) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001100) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001100) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001100) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001100) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001100) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001100) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001100) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001100) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001100) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001100) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001100) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001100) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001100) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001100) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001100) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001100) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001100) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001100) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001100) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001100) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001100) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001100) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001100) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001100) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001100) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001100) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001100) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001100) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001100) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001100) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001100) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001100) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001100) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001100) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001100) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001100) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001100) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001100) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001100) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001100) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001100) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001100) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001100) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001100) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001100) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001100) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001100) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001100) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001100) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001100) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001100) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001100) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001100) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001100) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001100) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001100) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001100) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001100) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001100) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001100) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001100) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001100) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001100) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001100) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001100) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001100) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001100) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001100) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001100) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001100) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001100) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001100) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001100) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001100) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001100) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001100) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001100) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001100) ? sw_input_81 :           
                    7'bzzzzzzz; 
assign sw_output_158 =(control_signal[1] == 1) ? stationary_signal_77:
                    
                     (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b1001101) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001101) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001101) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001101) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001101) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001101) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001101) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001101) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001101) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001101) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001101) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001101) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001101) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001101) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001101) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001101) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001101) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001101) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001101) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001101) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001101) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001101) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001101) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001101) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001101) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001101) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001101) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001101) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001101) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001101) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001101) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001101) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001101) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001101) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001101) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001101) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001101) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001101) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001101) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001101) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001101) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001101) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001101) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001101) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001101) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001101) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001101) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001101) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001101) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001101) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001101) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001101) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001101) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001101) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001101) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001101) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001101) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001101) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001101) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001101) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001101) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001101) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001101) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001101) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001101) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001101) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001101) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001101) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001101) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001101) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001101) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001101) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001101) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001101) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001101) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001101) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001101) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001101) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001101) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001101) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001101) ? sw_input_81 :            
                    7'bzzzzzzz; 
 assign sw_output_159 =(control_signal[1] == 1) ? stationary_signal_78:
                    
                     (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :
                    
                     (control_signal[0] ==0&& index_1 == 7'b1001110) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001110) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001110) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001110) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001110) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001110) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001110) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001110) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001110) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001110) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001110) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001110) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001110) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001110) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001110) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001110) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001110) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001110) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001110) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001110) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001110) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001110) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001110) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001110) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001110) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001110) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001110) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001110) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001110) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001110) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001110) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001110) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001110) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001110) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001110) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001110) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001110) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001110) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001110) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001110) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001110) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001110) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001110) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001110) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001110) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001110) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001110) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001110) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001110) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001110) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001110) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001110) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001110) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001110) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001110) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001110) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001110) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001110) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001110) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001110) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001110) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001110) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001110) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001110) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001110) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001110) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001110) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001110) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001110) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001110) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001110) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001110) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001110) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001110) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001110) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001110) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001110) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001110) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001110) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001110) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001110) ? sw_input_81 :            
                    7'bzzzzzzz; 
assign sw_output_160 =(control_signal[1] == 1) ? stationary_signal_79:

                     (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b1001111) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1001111) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1001111) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1001111) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1001111) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1001111) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1001111) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1001111) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1001111) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1001111) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1001111) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1001111) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1001111) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1001111) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1001111) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1001111) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1001111) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1001111) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1001111) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1001111) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1001111) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1001111) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1001111) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1001111) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1001111) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1001111) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1001111) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1001111) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1001111) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1001111) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1001111) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1001111) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1001111) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1001111) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1001111) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1001111) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1001111) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1001111) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1001111) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1001111) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1001111) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1001111) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1001111) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1001111) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1001111) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1001111) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1001111) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1001111) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1001111) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1001111) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1001111) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1001111) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1001111) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1001111) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1001111) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1001111) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1001111) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1001111) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1001111) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1001111) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1001111) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1001111) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1001111) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1001111) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1001111) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1001111) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1001111) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1001111) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1001111) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1001111) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1001111) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1001111) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1001111) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1001111) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1001111) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1001111) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1001111) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1001111) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1001111) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1001111) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1001111) ? sw_input_81 :            
                    7'bzzzzzzz; 
assign sw_output_161 =(control_signal[1] == 1) ? stationary_signal_80:

                     (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b1010000) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1010000) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1010000) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1010000) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1010000) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1010000) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1010000) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1010000) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1010000) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1010000) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1010000) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1010000) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1010000) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1010000) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1010000) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1010000) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1010000) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1010000) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1010000) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1010000) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1010000) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1010000) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1010000) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1010000) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1010000) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1010000) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1010000) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1010000) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1010000) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1010000) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1010000) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1010000) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1010000) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1010000) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1010000) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1010000) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1010000) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1010000) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1010000) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1010000) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1010000) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1010000) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1010000) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1010000) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1010000) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1010000) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1010000) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1010000) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1010000) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1010000) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1010000) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1010000) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1010000) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1010000) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1010000) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1010000) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1010000) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1010000) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1010000) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1010000) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1010000) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1010000) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1010000) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1010000) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1010000) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1010000) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1010000) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1010000) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1010000) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1010000) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1010000) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1010000) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1010000) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1010000) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1010000) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1010000) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1010000) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1010000) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1010000) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1010000) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1010000) ? sw_input_81 :             
                    7'bzzzzzzz; 
assign sw_output_162 =(control_signal[1] == 1) ? stationary_signal_81:
                      (control_signal[0] ==1&& index_1 == 7'b0001001) ? sw_input_1 :
                      (control_signal[0] ==1&& index_2 == 7'b0001001) ? sw_input_2 : 
                      (control_signal[0] ==1&& index_3 == 7'b0001001) ? sw_input_3 : 
                      (control_signal[0] ==1&& index_4 == 7'b0001001) ? sw_input_4 : 
                      (control_signal[0] ==1&& index_5 == 7'b0001001) ? sw_input_5 : 
                      (control_signal[0] ==1&& index_6 == 7'b0001001) ? sw_input_6 : 
                      (control_signal[0] ==1&& index_7 == 7'b0001001) ? sw_input_7 : 
                      (control_signal[0] ==1&& index_8 == 7'b0001001) ? sw_input_8 :
                      (control_signal[0] ==1&& index_9 == 7'b0001001) ? sw_input_9 :
                    
                    (control_signal[0] ==0&& index_1 == 7'b1010001) ? sw_input_1 : 
                    (control_signal[0] ==0&& index_2 == 7'b1010001) ? sw_input_2 : 
                    (control_signal[0] ==0&& index_3 == 7'b1010001) ? sw_input_3 : 
                    (control_signal[0] ==0&& index_4 == 7'b1010001) ? sw_input_4 : 
                    (control_signal[0] ==0&& index_5 == 7'b1010001) ? sw_input_5 : 
                    (control_signal[0] ==0&& index_6 == 7'b1010001) ? sw_input_6 : 
                    (control_signal[0] ==0&& index_7 == 7'b1010001) ? sw_input_7 : 
                    (control_signal[0] ==0&& index_8 == 7'b1010001) ? sw_input_8 :              
                    (control_signal[0] ==0&& index_9 == 7'b1010001) ? sw_input_9 : 
                    (control_signal[0] ==0&& index_10 == 7'b1010001) ? sw_input_10 : 
                    (control_signal[0] ==0&& index_11 == 7'b1010001) ? sw_input_11 : 
                    (control_signal[0] ==0&& index_12 == 7'b1010001) ? sw_input_12 : 
                    (control_signal[0] ==0&& index_13 == 7'b1010001) ? sw_input_13 : 
                    (control_signal[0] ==0&& index_14 == 7'b1010001) ? sw_input_14 : 
                    (control_signal[0] ==0&& index_15 == 7'b1010001) ? sw_input_15 : 
                    (control_signal[0] ==0&& index_16 == 7'b1010001) ? sw_input_16 : 
                    (control_signal[0] ==0&& index_17 == 7'b1010001) ? sw_input_17: 
                    (control_signal[0] ==0&& index_18 == 7'b1010001) ? sw_input_18 : 
                    (control_signal[0] ==0&& index_19 == 7'b1010001) ? sw_input_19 : 
                    (control_signal[0] ==0&& index_20 == 7'b1010001) ? sw_input_20 : 
                    (control_signal[0] ==0&& index_21 == 7'b1010001) ? sw_input_21 : 
                    (control_signal[0] ==0&& index_22 == 7'b1010001) ? sw_input_22 : 
                    (control_signal[0] ==0&& index_23 == 7'b1010001) ? sw_input_23 : 
                    (control_signal[0] ==0&& index_24 == 7'b1010001) ? sw_input_24 : 
                    (control_signal[0] ==0&& index_25 == 7'b1010001) ? sw_input_25 : 
                    (control_signal[0] ==0&& index_26 == 7'b1010001) ? sw_input_26 : 
                    (control_signal[0] ==0&& index_27 == 7'b1010001) ? sw_input_27 : 
                    (control_signal[0] ==0&& index_28 == 7'b1010001) ? sw_input_28 : 
                    (control_signal[0] ==0&& index_29 == 7'b1010001) ? sw_input_29 : 
                    (control_signal[0] ==0&& index_30 == 7'b1010001) ? sw_input_30 : 
                    (control_signal[0] ==0&& index_31 == 7'b1010001) ? sw_input_31 : 
                    (control_signal[0] ==0&& index_32 == 7'b1010001) ? sw_input_32 : 
                    (control_signal[0] ==0&& index_33 == 7'b1010001) ? sw_input_33 : 
                    (control_signal[0] ==0&& index_34 == 7'b1010001) ? sw_input_34 : 
                    (control_signal[0] ==0&& index_35 == 7'b1010001) ? sw_input_35 : 
                    (control_signal[0] ==0&& index_36 == 7'b1010001) ? sw_input_36 : 
                    (control_signal[0] ==0&& index_37 == 7'b1010001) ? sw_input_37 : 
                    (control_signal[0] ==0&& index_38 == 7'b1010001) ? sw_input_38 : 
                    (control_signal[0] ==0&& index_39 == 7'b1010001) ? sw_input_39 : 
                    (control_signal[0] ==0&& index_40 == 7'b1010001) ? sw_input_40 : 
                    (control_signal[0] ==0&& index_41 == 7'b1010001) ? sw_input_41 : 
                    (control_signal[0] ==0&& index_42 == 7'b1010001) ? sw_input_42 : 
                    (control_signal[0] ==0&& index_43 == 7'b1010001) ? sw_input_43 : 
                    (control_signal[0] ==0&& index_44 == 7'b1010001) ? sw_input_44 : 
                    (control_signal[0] ==0&& index_45 == 7'b1010001) ? sw_input_45 : 
                    (control_signal[0] ==0&& index_46 == 7'b1010001) ? sw_input_46 : 
                    (control_signal[0] ==0&& index_47 == 7'b1010001) ? sw_input_47 : 
                    (control_signal[0] ==0&& index_48 == 7'b1010001) ? sw_input_48 : 
                    (control_signal[0] ==0&& index_49 == 7'b1010001) ? sw_input_49 : 
                    (control_signal[0] ==0&& index_50 == 7'b1010001) ? sw_input_50 : 
                    (control_signal[0] ==0&& index_51 == 7'b1010001) ? sw_input_51 : 
                    (control_signal[0] ==0&& index_52 == 7'b1010001) ? sw_input_52 : 
                    (control_signal[0] ==0&& index_53 == 7'b1010001) ? sw_input_53 : 
                    (control_signal[0] ==0&& index_54 == 7'b1010001) ? sw_input_54 : 
                    (control_signal[0] ==0&& index_55 == 7'b1010001) ? sw_input_55 : 
                    (control_signal[0] ==0&& index_56 == 7'b1010001) ? sw_input_56 : 
                    (control_signal[0] ==0&& index_57 == 7'b1010001) ? sw_input_57 : 
                    (control_signal[0] ==0&& index_58 == 7'b1010001) ? sw_input_58 : 
                    (control_signal[0] ==0&& index_59 == 7'b1010001) ? sw_input_59 : 
                    (control_signal[0] ==0&& index_60 == 7'b1010001) ? sw_input_60 : 
                    (control_signal[0] ==0&& index_61 == 7'b1010001) ? sw_input_61 : 
                    (control_signal[0] ==0&& index_62 == 7'b1010001) ? sw_input_62 : 
                    (control_signal[0] ==0&& index_63 == 7'b1010001) ? sw_input_63 : 
                    (control_signal[0] ==0&& index_64 == 7'b1010001) ? sw_input_64 : 
                    (control_signal[0] ==0&& index_65 == 7'b1010001) ? sw_input_65 : 
                    (control_signal[0] ==0&& index_66 == 7'b1010001) ? sw_input_66 : 
                    (control_signal[0] ==0&& index_67 == 7'b1010001) ? sw_input_67 : 
                    (control_signal[0] ==0&& index_68 == 7'b1010001) ? sw_input_68 : 
                    (control_signal[0] ==0&& index_69 == 7'b1010001) ? sw_input_69 : 
                    (control_signal[0] ==0&& index_70 == 7'b1010001) ? sw_input_70 : 
                    (control_signal[0] ==0&& index_71 == 7'b1010001) ? sw_input_71 : 
                    (control_signal[0] ==0&& index_72 == 7'b1010001) ? sw_input_72 : 
                    (control_signal[0] ==0&& index_73 == 7'b1010001) ? sw_input_73 : 
                    (control_signal[0] ==0&& index_74 == 7'b1010001) ? sw_input_74 : 
                    (control_signal[0] ==0&& index_75 == 7'b1010001) ? sw_input_75 : 
                    (control_signal[0] ==0&& index_76 == 7'b1010001) ? sw_input_76 : 
                    (control_signal[0] ==0&& index_77 == 7'b1010001) ? sw_input_77 : 
                    (control_signal[0] ==0&& index_78 == 7'b1010001) ? sw_input_78 :  
                    (control_signal[0] ==0&& index_79 == 7'b1010001) ? sw_input_79 : 
                    (control_signal[0] ==0&& index_80 == 7'b1010001) ? sw_input_80 : 
                    (control_signal[0] ==0&& index_81 == 7'b1010001) ? sw_input_81 :
                                
                    7'bzzzzzzz; 
endmodule

