`timescale 10ns / 1ns



module tb_npu#(parameter WIDTH =4,INPUT_WIDTH = 9, INPUT_HEIGHT = 9,KERNEL_SIZE = 3,WEIGHT_HEIGHT = 3,WEIGHT_WIDTH = 3,PADDING_SIZE=0,STRIDE=1, batch_size = ((((((INPUT_HEIGHT-KERNEL_SIZE+(2*PADDING_SIZE)+1)/STRIDE))*(((INPUT_WIDTH-KERNEL_SIZE+(2*PADDING_SIZE)+1)/STRIDE))*9)-1)/81));
reg clk;
reg reset;
reg [31:0] axi_input_data;         
reg [31:0]axi_input_handshake;                     
reg [31:0] control_signal; 
wire [31:0] axi_output_data;
wire [31:0] axi_output_handshake;

      

npu inst_npu(                           //npu instantiation
.clk(clk),
.reset(reset),
.axi_input_data(axi_input_data),
.axi_input_handshake(axi_input_handshake),
.control_signal(control_signal),
.axi_output_data(axi_output_data),
.axi_output_handshake(axi_output_handshake)
    );
    
always begin                        //clock generation
    #5 clk = ~clk;
end
  
initial begin
    clk = 1;                
    reset = 1;
    
    #10
    
 // Testcase1 = Weight Stationary Unicast ,WIDTH =4,INPUT_WIDTH = 9, INPUT_HEIGHT = 9,KERNEL_SIZE = 3,WEIGHT_HEIGHT = 3,WEIGHT_WIDTH = 3,PADDING=0,STRIDE=1
 // ATTENTION : parameter declaration in all modules need to be changed when testing a new kind of stationary data flow
 // Testcase description : Testing weight stationary with Input size =9*9
 /*
 reset = 0;
control_signal =2'b00; 
axi_input_valid=1'b1;               
axi_input_ready=1'b1;

//inputs

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


#20;


//weights


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

#30;

//indexes
axi_input_data = 32'h1;   #10;
axi_input_data = 32'h2;   #10;
axi_input_data = 32'h3;   #10;
axi_input_data = 32'h4;   #10;
axi_input_data = 32'h5;   #10;
axi_input_data = 32'h6;   #10;
axi_input_data = 32'h7;   #10;
axi_input_data = 32'h8;   #10;
axi_input_data = 32'h9;   #10;
axi_input_data = 32'hA;   #10;
axi_input_data = 32'hB;   #10;
axi_input_data = 32'hC;   #10;
axi_input_data = 32'hD;   #10;
axi_input_data = 32'hE;   #10;
axi_input_data = 32'hF;   #10;
axi_input_data = 32'h10;  #10;
axi_input_data = 32'h11;  #10;
axi_input_data = 32'h12;  #10;
axi_input_data = 32'h13;  #10;
axi_input_data = 32'h14;  #10;
axi_input_data = 32'h15;  #10;
axi_input_data = 32'h16;  #10;
axi_input_data = 32'h17;  #10;
axi_input_data = 32'h18;  #10;
axi_input_data = 32'h19;  #10;
axi_input_data = 32'h1A;  #10;
axi_input_data = 32'h1B;  #10;
axi_input_data = 32'h1C;  #10;
axi_input_data = 32'h1D;  #10;
axi_input_data = 32'h1E;  #10;
axi_input_data = 32'h1F;  #10;
axi_input_data = 32'h20;  #10;
axi_input_data = 32'h21;  #10;
axi_input_data = 32'h22;  #10;
axi_input_data = 32'h23;  #10;
axi_input_data = 32'h24;  #10;
axi_input_data = 32'h25;  #10;
axi_input_data = 32'h26;  #10;
axi_input_data = 32'h27;  #10;
axi_input_data = 32'h28;  #10;
axi_input_data = 32'h29;  #10;
axi_input_data = 32'h2A;  #10;
axi_input_data = 32'h2B;  #10;
axi_input_data = 32'h2C;  #10;
axi_input_data = 32'h2D;  #10;
axi_input_data = 32'h2E;  #10;
axi_input_data = 32'h2F;  #10;
axi_input_data = 32'h30;  #10;
axi_input_data = 32'h31;  #10;
axi_input_data = 32'h32;  #10;
axi_input_data = 32'h33;  #10;
axi_input_data = 32'h34;  #10;
axi_input_data = 32'h35;  #10;
axi_input_data = 32'h36;  #10;
axi_input_data = 32'h37;  #10;
axi_input_data = 32'h38;  #10;
axi_input_data = 32'h39;  #10;
axi_input_data = 32'h3A;  #10;
axi_input_data = 32'h3B;  #10;
axi_input_data = 32'h3C;  #10;
axi_input_data = 32'h3D;  #10;
axi_input_data = 32'h3E;  #10;
axi_input_data = 32'h3F;  #10;
axi_input_data = 32'h40;  #10;
axi_input_data = 32'h41;  #10;
axi_input_data = 32'h42;  #10;
axi_input_data = 32'h43;  #10;
axi_input_data = 32'h44;  #10;
axi_input_data = 32'h45;  #10;
axi_input_data = 32'h46;  #10;
axi_input_data = 32'h47;  #10;
axi_input_data = 32'h48;  #10;
axi_input_data = 32'h49;  #10;
axi_input_data = 32'h4A;  #10;
axi_input_data = 32'h4B;  #10;
axi_input_data = 32'h4C;  #10;
axi_input_data = 32'h4D;  #10;
axi_input_data = 32'h4E;  #10;
axi_input_data = 32'h4F;  #10;
axi_input_data = 32'h50;  #10;
axi_input_data = 32'h51;  #10; */

// Testcase2 = Input Stationary Unicast ,WIDTH =4,INPUT_WIDTH = 9, INPUT_HEIGHT = 9,KERNEL_SIZE = 3,WEIGHT_HEIGHT = 21,WEIGHT_WIDTH = 21,PADDING=0,STRIDE=1
 // ATTENTION : parameter declaration in all modules need to be changed when testing a new kind of stationary data flow
  // Testcase description : Testing input stationary with Input size =9*9
 // the size of weight matrix should be equal to number of coefficients required=Here in  this case  7*7*9 =441
/*reset = 0;
control_signal =2'b10; 
axi_input_valid=1'b1;               
axi_input_ready=1'b1;

//inputs

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


#20;


//weights


axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;


//



axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;


//weights


axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;



#30;

//indexes
axi_input_data = 32'h1;   #10;
axi_input_data = 32'h2;   #10;
axi_input_data = 32'h3;   #10;
axi_input_data = 32'h4;   #10;
axi_input_data = 32'h5;   #10;
axi_input_data = 32'h6;   #10;
axi_input_data = 32'h7;   #10;
axi_input_data = 32'h8;   #10;
axi_input_data = 32'h9;   #10;
axi_input_data = 32'hA;   #10;
axi_input_data = 32'hB;   #10;
axi_input_data = 32'hC;   #10;
axi_input_data = 32'hD;   #10;
axi_input_data = 32'hE;   #10;
axi_input_data = 32'hF;   #10;
axi_input_data = 32'h10;  #10;
axi_input_data = 32'h11;  #10;
axi_input_data = 32'h12;  #10;
axi_input_data = 32'h13;  #10;
axi_input_data = 32'h14;  #10;
axi_input_data = 32'h15;  #10;
axi_input_data = 32'h16;  #10;
axi_input_data = 32'h17;  #10;
axi_input_data = 32'h18;  #10;
axi_input_data = 32'h19;  #10;
axi_input_data = 32'h1A;  #10;
axi_input_data = 32'h1B;  #10;
axi_input_data = 32'h1C;  #10;
axi_input_data = 32'h1D;  #10;
axi_input_data = 32'h1E;  #10;
axi_input_data = 32'h1F;  #10;
axi_input_data = 32'h20;  #10;
axi_input_data = 32'h21;  #10;
axi_input_data = 32'h22;  #10;
axi_input_data = 32'h23;  #10;
axi_input_data = 32'h24;  #10;
axi_input_data = 32'h25;  #10;
axi_input_data = 32'h26;  #10;
axi_input_data = 32'h27;  #10;
axi_input_data = 32'h28;  #10;
axi_input_data = 32'h29;  #10;
axi_input_data = 32'h2A;  #10;
axi_input_data = 32'h2B;  #10;
axi_input_data = 32'h2C;  #10;
axi_input_data = 32'h2D;  #10;
axi_input_data = 32'h2E;  #10;
axi_input_data = 32'h2F;  #10;
axi_input_data = 32'h30;  #10;
axi_input_data = 32'h31;  #10;
axi_input_data = 32'h32;  #10;
axi_input_data = 32'h33;  #10;
axi_input_data = 32'h34;  #10;
axi_input_data = 32'h35;  #10;
axi_input_data = 32'h36;  #10;
axi_input_data = 32'h37;  #10;
axi_input_data = 32'h38;  #10;
axi_input_data = 32'h39;  #10;
axi_input_data = 32'h3A;  #10;
axi_input_data = 32'h3B;  #10;
axi_input_data = 32'h3C;  #10;
axi_input_data = 32'h3D;  #10;
axi_input_data = 32'h3E;  #10;
axi_input_data = 32'h3F;  #10;
axi_input_data = 32'h40;  #10;
axi_input_data = 32'h41;  #10;
axi_input_data = 32'h42;  #10;
axi_input_data = 32'h43;  #10;
axi_input_data = 32'h44;  #10;
axi_input_data = 32'h45;  #10;
axi_input_data = 32'h46;  #10;
axi_input_data = 32'h47;  #10;
axi_input_data = 32'h48;  #10;
axi_input_data = 32'h49;  #10;
axi_input_data = 32'h4A;  #10;
axi_input_data = 32'h4B;  #10;
axi_input_data = 32'h4C;  #10;
axi_input_data = 32'h4D;  #10;
axi_input_data = 32'h4E;  #10;
axi_input_data = 32'h4F;  #10;
axi_input_data = 32'h50;  #10;
axi_input_data = 32'h51;  #10;*/


// Testcase3 = Input Stationary Unicast ,WIDTH =4,INPUT_WIDTH = 15, INPUT_HEIGHT = 15,KERNEL_SIZE = 3,WEIGHT_HEIGHT = 39,WEIGHT_WIDTH = 39,PADDING=0,STRIDE=1
// Testcase description : Testing input stationary with Input size =15*15
 // ATTENTION : parameter declaration in all modules need to be changed when testing a new kind of stationary data flow
 // the size of weight matrix should be equal to number of coefficients required=Here in  this case  7*7*9 =441

/*reset = 0;
control_signal =2'b10; 
axi_input_valid=1'b1;               
axi_input_ready=1'b1;

//inputs

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;


#20;


//weights


axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;


//weights


axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;


//weights


axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;


//weights


axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;


//weights


axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;


//weights


axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;


//weights


axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;


//weights


axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;


//weights


axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;






#30;

//indexes
axi_input_data = 32'h1;   #10;
axi_input_data = 32'h2;   #10;
axi_input_data = 32'h3;   #10;
axi_input_data = 32'h4;   #10;
axi_input_data = 32'h5;   #10;
axi_input_data = 32'h6;   #10;
axi_input_data = 32'h7;   #10;
axi_input_data = 32'h8;   #10;
axi_input_data = 32'h9;   #10;
axi_input_data = 32'hA;   #10;
axi_input_data = 32'hB;   #10;
axi_input_data = 32'hC;   #10;
axi_input_data = 32'hD;   #10;
axi_input_data = 32'hE;   #10;
axi_input_data = 32'hF;   #10;
axi_input_data = 32'h10;  #10;
axi_input_data = 32'h11;  #10;
axi_input_data = 32'h12;  #10;
axi_input_data = 32'h13;  #10;
axi_input_data = 32'h14;  #10;
axi_input_data = 32'h15;  #10;
axi_input_data = 32'h16;  #10;
axi_input_data = 32'h17;  #10;
axi_input_data = 32'h18;  #10;
axi_input_data = 32'h19;  #10;
axi_input_data = 32'h1A;  #10;
axi_input_data = 32'h1B;  #10;
axi_input_data = 32'h1C;  #10;
axi_input_data = 32'h1D;  #10;
axi_input_data = 32'h1E;  #10;
axi_input_data = 32'h1F;  #10;
axi_input_data = 32'h20;  #10;
axi_input_data = 32'h21;  #10;
axi_input_data = 32'h22;  #10;
axi_input_data = 32'h23;  #10;
axi_input_data = 32'h24;  #10;
axi_input_data = 32'h25;  #10;
axi_input_data = 32'h26;  #10;
axi_input_data = 32'h27;  #10;
axi_input_data = 32'h28;  #10;
axi_input_data = 32'h29;  #10;
axi_input_data = 32'h2A;  #10;
axi_input_data = 32'h2B;  #10;
axi_input_data = 32'h2C;  #10;
axi_input_data = 32'h2D;  #10;
axi_input_data = 32'h2E;  #10;
axi_input_data = 32'h2F;  #10;
axi_input_data = 32'h30;  #10;
axi_input_data = 32'h31;  #10;
axi_input_data = 32'h32;  #10;
axi_input_data = 32'h33;  #10;
axi_input_data = 32'h34;  #10;
axi_input_data = 32'h35;  #10;
axi_input_data = 32'h36;  #10;
axi_input_data = 32'h37;  #10;
axi_input_data = 32'h38;  #10;
axi_input_data = 32'h39;  #10;
axi_input_data = 32'h3A;  #10;
axi_input_data = 32'h3B;  #10;
axi_input_data = 32'h3C;  #10;
axi_input_data = 32'h3D;  #10;
axi_input_data = 32'h3E;  #10;
axi_input_data = 32'h3F;  #10;
axi_input_data = 32'h40;  #10;
axi_input_data = 32'h41;  #10;
axi_input_data = 32'h42;  #10;
axi_input_data = 32'h43;  #10;
axi_input_data = 32'h44;  #10;
axi_input_data = 32'h45;  #10;
axi_input_data = 32'h46;  #10;
axi_input_data = 32'h47;  #10;
axi_input_data = 32'h48;  #10;
axi_input_data = 32'h49;  #10;
axi_input_data = 32'h4A;  #10;
axi_input_data = 32'h4B;  #10;
axi_input_data = 32'h4C;  #10;
axi_input_data = 32'h4D;  #10;
axi_input_data = 32'h4E;  #10;
axi_input_data = 32'h4F;  #10;
axi_input_data = 32'h50;  #10;
axi_input_data = 32'h51;  #10;*/



// Testcase4 = Weight Stationary Unicast ,WIDTH =4,INPUT_WIDTH = 15, INPUT_HEIGHT = 15,KERNEL_SIZE = 3,WEIGHT_HEIGHT = 9,WEIGHT_WIDTH = 9,PADDING=0,STRIDE=1
// Testcase description : Testing Weight stationary with Input size =15*15
 // ATTENTION : parameter declaration in all modules need to be changed when testing a new kind of stationary data flow
 /*
reset = 0;
control_signal =2'b00; 
axi_input_valid=1'b1;               
axi_input_ready=1'b1;

//inputs

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;


#20;

//weights


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;






#30;

//indexes
axi_input_data = 32'h1;   #10;
axi_input_data = 32'h2;   #10;
axi_input_data = 32'h3;   #10;
axi_input_data = 32'h4;   #10;
axi_input_data = 32'h5;   #10;
axi_input_data = 32'h6;   #10;
axi_input_data = 32'h7;   #10;
axi_input_data = 32'h8;   #10;
axi_input_data = 32'h9;   #10;
axi_input_data = 32'hA;   #10;
axi_input_data = 32'hB;   #10;
axi_input_data = 32'hC;   #10;
axi_input_data = 32'hD;   #10;
axi_input_data = 32'hE;   #10;
axi_input_data = 32'hF;   #10;
axi_input_data = 32'h10;  #10;
axi_input_data = 32'h11;  #10;
axi_input_data = 32'h12;  #10;
axi_input_data = 32'h13;  #10;
axi_input_data = 32'h14;  #10;
axi_input_data = 32'h15;  #10;
axi_input_data = 32'h16;  #10;
axi_input_data = 32'h17;  #10;
axi_input_data = 32'h18;  #10;
axi_input_data = 32'h19;  #10;
axi_input_data = 32'h1A;  #10;
axi_input_data = 32'h1B;  #10;
axi_input_data = 32'h1C;  #10;
axi_input_data = 32'h1D;  #10;
axi_input_data = 32'h1E;  #10;
axi_input_data = 32'h1F;  #10;
axi_input_data = 32'h20;  #10;
axi_input_data = 32'h21;  #10;
axi_input_data = 32'h22;  #10;
axi_input_data = 32'h23;  #10;
axi_input_data = 32'h24;  #10;
axi_input_data = 32'h25;  #10;
axi_input_data = 32'h26;  #10;
axi_input_data = 32'h27;  #10;
axi_input_data = 32'h28;  #10;
axi_input_data = 32'h29;  #10;
axi_input_data = 32'h2A;  #10;
axi_input_data = 32'h2B;  #10;
axi_input_data = 32'h2C;  #10;
axi_input_data = 32'h2D;  #10;
axi_input_data = 32'h2E;  #10;
axi_input_data = 32'h2F;  #10;
axi_input_data = 32'h30;  #10;
axi_input_data = 32'h31;  #10;
axi_input_data = 32'h32;  #10;
axi_input_data = 32'h33;  #10;
axi_input_data = 32'h34;  #10;
axi_input_data = 32'h35;  #10;
axi_input_data = 32'h36;  #10;
axi_input_data = 32'h37;  #10;
axi_input_data = 32'h38;  #10;
axi_input_data = 32'h39;  #10;
axi_input_data = 32'h3A;  #10;
axi_input_data = 32'h3B;  #10;
axi_input_data = 32'h3C;  #10;
axi_input_data = 32'h3D;  #10;
axi_input_data = 32'h3E;  #10;
axi_input_data = 32'h3F;  #10;
axi_input_data = 32'h40;  #10;
axi_input_data = 32'h41;  #10;
axi_input_data = 32'h42;  #10;
axi_input_data = 32'h43;  #10;
axi_input_data = 32'h44;  #10;
axi_input_data = 32'h45;  #10;
axi_input_data = 32'h46;  #10;
axi_input_data = 32'h47;  #10;
axi_input_data = 32'h48;  #10;
axi_input_data = 32'h49;  #10;
axi_input_data = 32'h4A;  #10;
axi_input_data = 32'h4B;  #10;
axi_input_data = 32'h4C;  #10;
axi_input_data = 32'h4D;  #10;
axi_input_data = 32'h4E;  #10;
axi_input_data = 32'h4F;  #10;
axi_input_data = 32'h50;  #10;
axi_input_data = 32'h51;  #10;
*/

 // Testcase5 = Weight Stationary Unicast ,WIDTH =8,INPUT_WIDTH = 9, INPUT_HEIGHT = 9,KERNEL_SIZE = 3,WEIGHT_HEIGHT = 3,WEIGHT_WIDTH = 3,PADDING=0,STRIDE=1
 // ATTENTION : parameter declaration in all modules need to be changed when testing a new kind of stationary data flow
 // Testcase description : Testing  bit width=8 for Weight stationary
 /*
reset = 0;
control_signal =2'b00; 
axi_input_valid=1'b1;               
axi_input_ready=1'b1;

//inputs

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


#20;


//weights


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

#30;

//indexes
axi_input_data = 32'h1;   #10;
axi_input_data = 32'h2;   #10;
axi_input_data = 32'h3;   #10;
axi_input_data = 32'h4;   #10;
axi_input_data = 32'h5;   #10;
axi_input_data = 32'h6;   #10;
axi_input_data = 32'h7;   #10;
axi_input_data = 32'h8;   #10;
axi_input_data = 32'h9;   #10;
axi_input_data = 32'hA;   #10;
axi_input_data = 32'hB;   #10;
axi_input_data = 32'hC;   #10;
axi_input_data = 32'hD;   #10;
axi_input_data = 32'hE;   #10;
axi_input_data = 32'hF;   #10;
axi_input_data = 32'h10;  #10;
axi_input_data = 32'h11;  #10;
axi_input_data = 32'h12;  #10;
axi_input_data = 32'h13;  #10;
axi_input_data = 32'h14;  #10;
axi_input_data = 32'h15;  #10;
axi_input_data = 32'h16;  #10;
axi_input_data = 32'h17;  #10;
axi_input_data = 32'h18;  #10;
axi_input_data = 32'h19;  #10;
axi_input_data = 32'h1A;  #10;
axi_input_data = 32'h1B;  #10;
axi_input_data = 32'h1C;  #10;
axi_input_data = 32'h1D;  #10;
axi_input_data = 32'h1E;  #10;
axi_input_data = 32'h1F;  #10;
axi_input_data = 32'h20;  #10;
axi_input_data = 32'h21;  #10;
axi_input_data = 32'h22;  #10;
axi_input_data = 32'h23;  #10;
axi_input_data = 32'h24;  #10;
axi_input_data = 32'h25;  #10;
axi_input_data = 32'h26;  #10;
axi_input_data = 32'h27;  #10;
axi_input_data = 32'h28;  #10;
axi_input_data = 32'h29;  #10;
axi_input_data = 32'h2A;  #10;
axi_input_data = 32'h2B;  #10;
axi_input_data = 32'h2C;  #10;
axi_input_data = 32'h2D;  #10;
axi_input_data = 32'h2E;  #10;
axi_input_data = 32'h2F;  #10;
axi_input_data = 32'h30;  #10;
axi_input_data = 32'h31;  #10;
axi_input_data = 32'h32;  #10;
axi_input_data = 32'h33;  #10;
axi_input_data = 32'h34;  #10;
axi_input_data = 32'h35;  #10;
axi_input_data = 32'h36;  #10;
axi_input_data = 32'h37;  #10;
axi_input_data = 32'h38;  #10;
axi_input_data = 32'h39;  #10;
axi_input_data = 32'h3A;  #10;
axi_input_data = 32'h3B;  #10;
axi_input_data = 32'h3C;  #10;
axi_input_data = 32'h3D;  #10;
axi_input_data = 32'h3E;  #10;
axi_input_data = 32'h3F;  #10;
axi_input_data = 32'h40;  #10;
axi_input_data = 32'h41;  #10;
axi_input_data = 32'h42;  #10;
axi_input_data = 32'h43;  #10;
axi_input_data = 32'h44;  #10;
axi_input_data = 32'h45;  #10;
axi_input_data = 32'h46;  #10;
axi_input_data = 32'h47;  #10;
axi_input_data = 32'h48;  #10;
axi_input_data = 32'h49;  #10;
axi_input_data = 32'h4A;  #10;
axi_input_data = 32'h4B;  #10;
axi_input_data = 32'h4C;  #10;
axi_input_data = 32'h4D;  #10;
axi_input_data = 32'h4E;  #10;
axi_input_data = 32'h4F;  #10;
axi_input_data = 32'h50;  #10;
axi_input_data = 32'h51;  #10; */

// Testcase6 = Weight Stationary Unicast ,WIDTH =8,INPUT_WIDTH = 5, INPUT_HEIGHT = 5,KERNEL_SIZE = 3,WEIGHT_HEIGHT = 3,WEIGHT_WIDTH = 3,PADDING=0,STRIDE=1
 // ATTENTION : parameter declaration in all modules need to be changed when testing a new kind of stationary data flow
 // Testcase description : Testing weight stationary with input size =5*5 and bit width =8
 
/*reset = 0;
control_signal =2'b00; 
axi_input_valid=1'b1;               
axi_input_ready=1'b1;

//inputs

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;





#20;


//weights


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

#30;

//indexes
axi_input_data = 32'h1;   #10;
axi_input_data = 32'h2;   #10;
axi_input_data = 32'h3;   #10;
axi_input_data = 32'h4;   #10;
axi_input_data = 32'h5;   #10;
axi_input_data = 32'h6;   #10;
axi_input_data = 32'h7;   #10;
axi_input_data = 32'h8;   #10;
axi_input_data = 32'h9;   #10;
axi_input_data = 32'hA;   #10;
axi_input_data = 32'hB;   #10;
axi_input_data = 32'hC;   #10;
axi_input_data = 32'hD;   #10;
axi_input_data = 32'hE;   #10;
axi_input_data = 32'hF;   #10;
axi_input_data = 32'h10;  #10;
axi_input_data = 32'h11;  #10;
axi_input_data = 32'h12;  #10;
axi_input_data = 32'h13;  #10;
axi_input_data = 32'h14;  #10;
axi_input_data = 32'h15;  #10;
axi_input_data = 32'h16;  #10;
axi_input_data = 32'h17;  #10;
axi_input_data = 32'h18;  #10;
axi_input_data = 32'h19;  #10;
axi_input_data = 32'h1A;  #10;
axi_input_data = 32'h1B;  #10;
axi_input_data = 32'h1C;  #10;
axi_input_data = 32'h1D;  #10;
axi_input_data = 32'h1E;  #10;
axi_input_data = 32'h1F;  #10;
axi_input_data = 32'h20;  #10;
axi_input_data = 32'h21;  #10;
axi_input_data = 32'h22;  #10;
axi_input_data = 32'h23;  #10;
axi_input_data = 32'h24;  #10;
axi_input_data = 32'h25;  #10;
axi_input_data = 32'h26;  #10;
axi_input_data = 32'h27;  #10;
axi_input_data = 32'h28;  #10;
axi_input_data = 32'h29;  #10;
axi_input_data = 32'h2A;  #10;
axi_input_data = 32'h2B;  #10;
axi_input_data = 32'h2C;  #10;
axi_input_data = 32'h2D;  #10;
axi_input_data = 32'h2E;  #10;
axi_input_data = 32'h2F;  #10;
axi_input_data = 32'h30;  #10;
axi_input_data = 32'h31;  #10;
axi_input_data = 32'h32;  #10;
axi_input_data = 32'h33;  #10;
axi_input_data = 32'h34;  #10;
axi_input_data = 32'h35;  #10;
axi_input_data = 32'h36;  #10;
axi_input_data = 32'h37;  #10;
axi_input_data = 32'h38;  #10;
axi_input_data = 32'h39;  #10;
axi_input_data = 32'h3A;  #10;
axi_input_data = 32'h3B;  #10;
axi_input_data = 32'h3C;  #10;
axi_input_data = 32'h3D;  #10;
axi_input_data = 32'h3E;  #10;
axi_input_data = 32'h3F;  #10;
axi_input_data = 32'h40;  #10;
axi_input_data = 32'h41;  #10;
axi_input_data = 32'h42;  #10;
axi_input_data = 32'h43;  #10;
axi_input_data = 32'h44;  #10;
axi_input_data = 32'h45;  #10;
axi_input_data = 32'h46;  #10;
axi_input_data = 32'h47;  #10;
axi_input_data = 32'h48;  #10;
axi_input_data = 32'h49;  #10;
axi_input_data = 32'h4A;  #10;
axi_input_data = 32'h4B;  #10;
axi_input_data = 32'h4C;  #10;
axi_input_data = 32'h4D;  #10;
axi_input_data = 32'h4E;  #10;
axi_input_data = 32'h4F;  #10;
axi_input_data = 32'h50;  #10;
axi_input_data = 32'h51;  #10;

*/


// Testcase7 = Weight Stationary Unicast ,WIDTH =4,INPUT_WIDTH = 64, INPUT_HEIGHT = 64,KERNEL_SIZE = 3,WEIGHT_HEIGHT = 3,WEIGHT_WIDTH = 3,PADDING=0,STRIDE=1
 // ATTENTION : parameter declaration in all modules need to be changed when testing a new kind of stationary data flow
 // Testcase description : Testing weight stationary with Input size =64*64
 /*
 reset = 0;
control_signal =2'b00; 
axi_input_valid=1'b1;               
axi_input_ready=1'b1;

//inputs

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;


#20;


//weights


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

#30;

//indexes
axi_input_data = 32'h1;   #10;
axi_input_data = 32'h2;   #10;
axi_input_data = 32'h3;   #10;
axi_input_data = 32'h4;   #10;
axi_input_data = 32'h5;   #10;
axi_input_data = 32'h6;   #10;
axi_input_data = 32'h7;   #10;
axi_input_data = 32'h8;   #10;
axi_input_data = 32'h9;   #10;
axi_input_data = 32'hA;   #10;
axi_input_data = 32'hB;   #10;
axi_input_data = 32'hC;   #10;
axi_input_data = 32'hD;   #10;
axi_input_data = 32'hE;   #10;
axi_input_data = 32'hF;   #10;
axi_input_data = 32'h10;  #10;
axi_input_data = 32'h11;  #10;
axi_input_data = 32'h12;  #10;
axi_input_data = 32'h13;  #10;
axi_input_data = 32'h14;  #10;
axi_input_data = 32'h15;  #10;
axi_input_data = 32'h16;  #10;
axi_input_data = 32'h17;  #10;
axi_input_data = 32'h18;  #10;
axi_input_data = 32'h19;  #10;
axi_input_data = 32'h1A;  #10;
axi_input_data = 32'h1B;  #10;
axi_input_data = 32'h1C;  #10;
axi_input_data = 32'h1D;  #10;
axi_input_data = 32'h1E;  #10;
axi_input_data = 32'h1F;  #10;
axi_input_data = 32'h20;  #10;
axi_input_data = 32'h21;  #10;
axi_input_data = 32'h22;  #10;
axi_input_data = 32'h23;  #10;
axi_input_data = 32'h24;  #10;
axi_input_data = 32'h25;  #10;
axi_input_data = 32'h26;  #10;
axi_input_data = 32'h27;  #10;
axi_input_data = 32'h28;  #10;
axi_input_data = 32'h29;  #10;
axi_input_data = 32'h2A;  #10;
axi_input_data = 32'h2B;  #10;
axi_input_data = 32'h2C;  #10;
axi_input_data = 32'h2D;  #10;
axi_input_data = 32'h2E;  #10;
axi_input_data = 32'h2F;  #10;
axi_input_data = 32'h30;  #10;
axi_input_data = 32'h31;  #10;
axi_input_data = 32'h32;  #10;
axi_input_data = 32'h33;  #10;
axi_input_data = 32'h34;  #10;
axi_input_data = 32'h35;  #10;
axi_input_data = 32'h36;  #10;
axi_input_data = 32'h37;  #10;
axi_input_data = 32'h38;  #10;
axi_input_data = 32'h39;  #10;
axi_input_data = 32'h3A;  #10;
axi_input_data = 32'h3B;  #10;
axi_input_data = 32'h3C;  #10;
axi_input_data = 32'h3D;  #10;
axi_input_data = 32'h3E;  #10;
axi_input_data = 32'h3F;  #10;
axi_input_data = 32'h40;  #10;
axi_input_data = 32'h41;  #10;
axi_input_data = 32'h42;  #10;
axi_input_data = 32'h43;  #10;
axi_input_data = 32'h44;  #10;
axi_input_data = 32'h45;  #10;
axi_input_data = 32'h46;  #10;
axi_input_data = 32'h47;  #10;
axi_input_data = 32'h48;  #10;
axi_input_data = 32'h49;  #10;
axi_input_data = 32'h4A;  #10;
axi_input_data = 32'h4B;  #10;
axi_input_data = 32'h4C;  #10;
axi_input_data = 32'h4D;  #10;
axi_input_data = 32'h4E;  #10;
axi_input_data = 32'h4F;  #10;
axi_input_data = 32'h50;  #10;
axi_input_data = 32'h51;  #10;
*/

// Testcase8 = Input Stationary Unicast ,WIDTH =4,INPUT_WIDTH = 7, INPUT_HEIGHT = 7,KERNEL_SIZE = 3,WEIGHT_HEIGHT = 21,WEIGHT_WIDTH = 21,PADDING=1,STRIDE=1
 // ATTENTION : parameter declaration in all modules need to be changed when testing a new kind of stationary data flow
  // Testcase description : Testing input stationary with Input size =7*7 with zero padding
/*
reset = 0;
control_signal =2'b10; 
axi_input_valid=1'b1;               
axi_input_ready=1'b1;

//inputs

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'hA;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'hD;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'hE;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'hA;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'hA;  #10;
axi_input_data = 32'hB;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;




#20;


//weights


axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h1;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;


//



axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;


//weights


axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h9;  #10;

//weights


axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h2;  #10;

axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h3;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;



#30;

//indexes
axi_input_data = 32'h1;   #10;
axi_input_data = 32'h2;   #10;
axi_input_data = 32'h3;   #10;
axi_input_data = 32'h4;   #10;
axi_input_data = 32'h5;   #10;
axi_input_data = 32'h6;   #10;
axi_input_data = 32'h7;   #10;
axi_input_data = 32'h8;   #10;
axi_input_data = 32'h9;   #10;
axi_input_data = 32'hA;   #10;
axi_input_data = 32'hB;   #10;
axi_input_data = 32'hC;   #10;
axi_input_data = 32'hD;   #10;
axi_input_data = 32'hE;   #10;
axi_input_data = 32'hF;   #10;
axi_input_data = 32'h10;  #10;
axi_input_data = 32'h11;  #10;
axi_input_data = 32'h12;  #10;
axi_input_data = 32'h13;  #10;
axi_input_data = 32'h14;  #10;
axi_input_data = 32'h15;  #10;
axi_input_data = 32'h16;  #10;
axi_input_data = 32'h17;  #10;
axi_input_data = 32'h18;  #10;
axi_input_data = 32'h19;  #10;
axi_input_data = 32'h1A;  #10;
axi_input_data = 32'h1B;  #10;
axi_input_data = 32'h1C;  #10;
axi_input_data = 32'h1D;  #10;
axi_input_data = 32'h1E;  #10;
axi_input_data = 32'h1F;  #10;
axi_input_data = 32'h20;  #10;
axi_input_data = 32'h21;  #10;
axi_input_data = 32'h22;  #10;
axi_input_data = 32'h23;  #10;
axi_input_data = 32'h24;  #10;
axi_input_data = 32'h25;  #10;
axi_input_data = 32'h26;  #10;
axi_input_data = 32'h27;  #10;
axi_input_data = 32'h28;  #10;
axi_input_data = 32'h29;  #10;
axi_input_data = 32'h2A;  #10;
axi_input_data = 32'h2B;  #10;
axi_input_data = 32'h2C;  #10;
axi_input_data = 32'h2D;  #10;
axi_input_data = 32'h2E;  #10;
axi_input_data = 32'h2F;  #10;
axi_input_data = 32'h30;  #10;
axi_input_data = 32'h31;  #10;
axi_input_data = 32'h32;  #10;
axi_input_data = 32'h33;  #10;
axi_input_data = 32'h34;  #10;
axi_input_data = 32'h35;  #10;
axi_input_data = 32'h36;  #10;
axi_input_data = 32'h37;  #10;
axi_input_data = 32'h38;  #10;
axi_input_data = 32'h39;  #10;
axi_input_data = 32'h3A;  #10;
axi_input_data = 32'h3B;  #10;
axi_input_data = 32'h3C;  #10;
axi_input_data = 32'h3D;  #10;
axi_input_data = 32'h3E;  #10;
axi_input_data = 32'h3F;  #10;
axi_input_data = 32'h40;  #10;
axi_input_data = 32'h41;  #10;
axi_input_data = 32'h42;  #10;
axi_input_data = 32'h43;  #10;
axi_input_data = 32'h44;  #10;
axi_input_data = 32'h45;  #10;
axi_input_data = 32'h46;  #10;
axi_input_data = 32'h47;  #10;
axi_input_data = 32'h48;  #10;
axi_input_data = 32'h49;  #10;
axi_input_data = 32'h4A;  #10;
axi_input_data = 32'h4B;  #10;
axi_input_data = 32'h4C;  #10;
axi_input_data = 32'h4D;  #10;
axi_input_data = 32'h4E;  #10;
axi_input_data = 32'h4F;  #10;
axi_input_data = 32'h50;  #10;
axi_input_data = 32'h51;  #10;  */

// Testcase9 = Weight Stationary Unicast ,WIDTH =8,INPUT_WIDTH = 32, INPUT_HEIGHT = 32,KERNEL_SIZE = 3,WEIGHT_HEIGHT = 3,WEIGHT_WIDTH = 3,PADDING=0,STRIDE=2
// Testcase description : Testing Weight stationary with Input size =32*32 and stride =2
 // ATTENTION : parameter declaration in all modules need to be changed when testing a new kind of stationary data flow
/*
reset = 0;
control_signal =2'b00; 
axi_input_valid=1'b1;               
axi_input_ready=1'b1;

//inputs

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'hC;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h15;  #10;

axi_input_data = 32'hC;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'hD;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h38;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'hD;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h48;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'hA;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h22;  #10;
axi_input_data = 32'hC;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h22;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h57;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5A;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h9;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'hA;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'hA;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h22;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10




#20;

//weights


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;






#30;

//indexes
axi_input_data = 32'h1;   #10;
axi_input_data = 32'h2;   #10;
axi_input_data = 32'h3;   #10;
axi_input_data = 32'h4;   #10;
axi_input_data = 32'h5;   #10;
axi_input_data = 32'h6;   #10;
axi_input_data = 32'h7;   #10;
axi_input_data = 32'h8;   #10;
axi_input_data = 32'h9;   #10;
axi_input_data = 32'hA;   #10;
axi_input_data = 32'hB;   #10;
axi_input_data = 32'hC;   #10;
axi_input_data = 32'hD;   #10;
axi_input_data = 32'hE;   #10;
axi_input_data = 32'hF;   #10;
axi_input_data = 32'h10;  #10;
axi_input_data = 32'h11;  #10;
axi_input_data = 32'h12;  #10;
axi_input_data = 32'h13;  #10;
axi_input_data = 32'h14;  #10;
axi_input_data = 32'h15;  #10;
axi_input_data = 32'h16;  #10;
axi_input_data = 32'h17;  #10;
axi_input_data = 32'h18;  #10;
axi_input_data = 32'h19;  #10;
axi_input_data = 32'h1A;  #10;
axi_input_data = 32'h1B;  #10;
axi_input_data = 32'h1C;  #10;
axi_input_data = 32'h1D;  #10;
axi_input_data = 32'h1E;  #10;
axi_input_data = 32'h1F;  #10;
axi_input_data = 32'h20;  #10;
axi_input_data = 32'h21;  #10;
axi_input_data = 32'h22;  #10;
axi_input_data = 32'h23;  #10;
axi_input_data = 32'h24;  #10;
axi_input_data = 32'h25;  #10;
axi_input_data = 32'h26;  #10;
axi_input_data = 32'h27;  #10;
axi_input_data = 32'h28;  #10;
axi_input_data = 32'h29;  #10;
axi_input_data = 32'h2A;  #10;
axi_input_data = 32'h2B;  #10;
axi_input_data = 32'h2C;  #10;
axi_input_data = 32'h2D;  #10;
axi_input_data = 32'h2E;  #10;
axi_input_data = 32'h2F;  #10;
axi_input_data = 32'h30;  #10;
axi_input_data = 32'h31;  #10;
axi_input_data = 32'h32;  #10;
axi_input_data = 32'h33;  #10;
axi_input_data = 32'h34;  #10;
axi_input_data = 32'h35;  #10;
axi_input_data = 32'h36;  #10;
axi_input_data = 32'h37;  #10;
axi_input_data = 32'h38;  #10;
axi_input_data = 32'h39;  #10;
axi_input_data = 32'h3A;  #10;
axi_input_data = 32'h3B;  #10;
axi_input_data = 32'h3C;  #10;
axi_input_data = 32'h3D;  #10;
axi_input_data = 32'h3E;  #10;
axi_input_data = 32'h3F;  #10;
axi_input_data = 32'h40;  #10;
axi_input_data = 32'h41;  #10;
axi_input_data = 32'h42;  #10;
axi_input_data = 32'h43;  #10;
axi_input_data = 32'h44;  #10;
axi_input_data = 32'h45;  #10;
axi_input_data = 32'h46;  #10;
axi_input_data = 32'h47;  #10;
axi_input_data = 32'h48;  #10;
axi_input_data = 32'h49;  #10;
axi_input_data = 32'h4A;  #10;
axi_input_data = 32'h4B;  #10;
axi_input_data = 32'h4C;  #10;
axi_input_data = 32'h4D;  #10;
axi_input_data = 32'h4E;  #10;
axi_input_data = 32'h4F;  #10;
axi_input_data = 32'h50;  #10;
axi_input_data = 32'h51;  #10;

*/
// Testcase11 = Final testcase to run on FPGA
//Weight Stationary Unicast ,WIDTH =4,INPUT_WIDTH = 9, INPUT_HEIGHT = 9,KERNEL_SIZE = 3,WEIGHT_HEIGHT = 3,WEIGHT_WIDTH = 3,PADDING=0,STRIDE=1
 // ATTENTION : parameter declaration in all modules need to be changed when testing a new kind of stationary data flow
 // Testcase description : Testing weight stationary with Input size =9*9
 
 reset = 0;
control_signal =32'b00; 
axi_input_handshake=32'd1;               


//inputs

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h0;  #10;

axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h4;  #10;

axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h5;  #10;

axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h6;  #10;

axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h7;  #10;

axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;
axi_input_data = 32'h8;  #10;


#20;


//weights


axi_input_data = 32'h0;  #10;
axi_input_data = 32'h1;  #10;
axi_input_data = 32'h2;  #10;
axi_input_data = 32'h3;  #10;
axi_input_data = 32'h4;  #10;
axi_input_data = 32'h5;  #10;
axi_input_data = 32'h6;  #10;
axi_input_data = 32'h7;  #10;
axi_input_data = 32'h8;  #10;

#30;

//indexes
axi_input_data = 32'h1;   #10;
axi_input_data = 32'h2;   #10;
axi_input_data = 32'h3;   #10;
axi_input_data = 32'h4;   #10;
axi_input_data = 32'h5;   #10;
axi_input_data = 32'h6;   #10;
axi_input_data = 32'h7;   #10;
axi_input_data = 32'h8;   #10;
axi_input_data = 32'h9;   #10;
axi_input_data = 32'hA;   #10;
axi_input_data = 32'hB;   #10;
axi_input_data = 32'hC;   #10;
axi_input_data = 32'hD;   #10;
axi_input_data = 32'hE;   #10;
axi_input_data = 32'hF;   #10;
axi_input_data = 32'h10;  #10;
axi_input_data = 32'h11;  #10;
axi_input_data = 32'h12;  #10;
axi_input_data = 32'h13;  #10;
axi_input_data = 32'h14;  #10;
axi_input_data = 32'h15;  #10;
axi_input_data = 32'h16;  #10;
axi_input_data = 32'h17;  #10;
axi_input_data = 32'h18;  #10;
axi_input_data = 32'h19;  #10;
axi_input_data = 32'h1A;  #10;
axi_input_data = 32'h1B;  #10;
axi_input_data = 32'h1C;  #10;
axi_input_data = 32'h1D;  #10;
axi_input_data = 32'h1E;  #10;
axi_input_data = 32'h1F;  #10;
axi_input_data = 32'h20;  #10;
axi_input_data = 32'h21;  #10;
axi_input_data = 32'h22;  #10;
axi_input_data = 32'h23;  #10;
axi_input_data = 32'h24;  #10;
axi_input_data = 32'h25;  #10;
axi_input_data = 32'h26;  #10;
axi_input_data = 32'h27;  #10;
axi_input_data = 32'h28;  #10;
axi_input_data = 32'h29;  #10;
axi_input_data = 32'h2A;  #10;
axi_input_data = 32'h2B;  #10;
axi_input_data = 32'h2C;  #10;
axi_input_data = 32'h2D;  #10;
axi_input_data = 32'h2E;  #10;
axi_input_data = 32'h2F;  #10;
axi_input_data = 32'h30;  #10;
axi_input_data = 32'h31;  #10;
axi_input_data = 32'h32;  #10;
axi_input_data = 32'h33;  #10;
axi_input_data = 32'h34;  #10;
axi_input_data = 32'h35;  #10;
axi_input_data = 32'h36;  #10;
axi_input_data = 32'h37;  #10;
axi_input_data = 32'h38;  #10;
axi_input_data = 32'h39;  #10;
axi_input_data = 32'h3A;  #10;
axi_input_data = 32'h3B;  #10;
axi_input_data = 32'h3C;  #10;
axi_input_data = 32'h3D;  #10;
axi_input_data = 32'h3E;  #10;
axi_input_data = 32'h3F;  #10;
axi_input_data = 32'h40;  #10;
axi_input_data = 32'h41;  #10;
axi_input_data = 32'h42;  #10;
axi_input_data = 32'h43;  #10;
axi_input_data = 32'h44;  #10;
axi_input_data = 32'h45;  #10;
axi_input_data = 32'h46;  #10;
axi_input_data = 32'h47;  #10;
axi_input_data = 32'h48;  #10;
axi_input_data = 32'h49;  #10;
axi_input_data = 32'h4A;  #10;
axi_input_data = 32'h4B;  #10;
axi_input_data = 32'h4C;  #10;
axi_input_data = 32'h4D;  #10;
axi_input_data = 32'h4E;  #10;
axi_input_data = 32'h4F;  #10;
axi_input_data = 32'h50;  #10;
axi_input_data = 32'h51;  #10;

#5000;
$finish;
end

endmodule

